`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Ronny Zarate Ferreto
// 
// Create Date: 26.09.2017 07:13:33
// Design Name: 
// Module Name: ROM_imagen_final
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ROM_imagen_final(
	input wire main_clk_i,
    input wire [8:0] address_i,
    output wire [0:639] data_o,
    output wire [9:0] W_o,
    output wire [8:0] H_o
    );
    
    //Registros
    reg [9:0] wREG; 
    reg [8:0] hREG; 
    reg [0:639] dataREG; 
    
    //ROM
    always @(posedge main_clk_i)
    begin
    hREG <= 480;
    wREG <= 640;
    case (address_i)
        
    0: dataREG =   640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000011111100011111000000000001111111111111000000001011111111111111111111111111111111111111111111010000000000000000000000000000000000000000000000000000000010111111000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    1: dataREG =   641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111010000000000000001111110111110000000000111111111111100000011111111111110110100001000000001010010101111111111111111100000000000000000000000000000000000000000000000000000011111111000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    2: dataREG =   641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000001111110011111010000001011111111100000111110111110101001000001000000000000000000000000000101111111111110100000000000000000000000000000000000000000000000000001111111000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    3: dataREG =   641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000111111111110000000011111111101101011011111010010000000000000000000000000000000000000100100000101111111111100000000000000000000000000000000000000000000000001011111110000000000000001110111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    5: dataREG =   641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011110110000000000001111111110110000001111011111101111111111010000000000000000000000001000000000000000000000000010000101011110111100000000000000000000000000000000000000000000000000111111100000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    6: dataREG =   641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111111000000000000111111111100000101111111101111101111000000000000000000000000000000000000000000000100000000000000000100011111110100000000000000000000000000000000000000000000000000111111000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    7: dataREG =   641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110110000000000111111111110000011011111111111111000000000000000000000000000000000000000000000000000000000000000000001000010111110110000100000000000000000000000000000000000000000010111111000000000101101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    9: dataREG =   641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101000010001011011111110001111111111111010100000000001000000000000000000000000000000000000000000000000000000000000100000100110111110111111110000000000000000000000000000000000000011101100000010111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    10: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001111110100000001111111111000010111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111111111010111100000000000000000000000000000000000000111110101011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    11: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000111111000000001111111101100011111110111010100001000000000000000000000000000000000000000000000000000000000000000000000000000000000001011101111111110100000000000000000000000000000001000101111011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    12: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111000000001111110000000111101011000111111111110000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100111111111111010000000000000000000000000000000000000111111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    13: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010000001111111000011011100000000111111111010000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000001111011111101010000100010000000000100000000000000001111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    14: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100100000111111000001111010000010111111100000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000011111111111101100010000010000000000000000000000000101101111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    15: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011110000000101111100111111100000011111101000000000000000000000000000000100010010010100100010000000000000000000010000000000000000000000000000000000000101111111111111100000000000000000000000000000000011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    16: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000011111110011111100000011111110010000000100001000000000001011001101101101010111101011010100010000100000000000000000000000000000000100000000000101111111111111100000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    17: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000111110101111100000011011000000000000011101111010000101111111111111111111111111111111111111110010001000000000000000000000000000000000000000011011111110111111000000000000000000000000000000000111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    18: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000111111111101000101111110000000001111111111111111111111111111111101111010101110111111111011111111110110010000000000000000000000000000000000000101111111111111111000000000000000000000000000000101111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    19: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001110010001011111111111000000111100000001011111111111111111111101001000000010000000010000000000001011011111111111110101000000000000000000000000000000000000111111111111110110000000000000000000000000010011011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    20: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110001111111101000011111000000101111101011101001010000000000000000000000010000000000000000000100000101111111111111100000000000000000000000100000000000111101111111111100000000000100010000000000000011111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    21: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101111111111000001111100000111110100000101000000000000000000000000000000000000000000000000000000000001011111111111101000000000100000000000000000010011110111111011111010000000000000000000000000001111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    22: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000111111100000111100000111101010000100001101101000010000000000000000000000000000000000000000000000000000001011111111110100000000000000000000000000001111111111111111001000000000000000000000000001111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    23: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110011101111001111111000000011100111101110000010111111110110000000000010000000000000000000000000000000000000000000000100101011111111010000000000000000000000000000111111011111111111010000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    24: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000010111100001111111011110000101111111111111100000000000000000000000000000000000000000000000001000000000000000100101111111110101000000000000000000000001011111111111111110000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    25: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011111111000001010100000111101111111111111110111101111110110000000000000000000000000000010000000000000000000000000000000000000011111111100100000000001000000000000101111010111111111100000000000000000000000001110111011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    26: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000010000011011111101101011111111111111011110111010000000000000000000000000000000000000000000000000000000000000000000111111111110100000000000000000000001011110111101011110100000000000000000000001111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    27: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000111111111110000000000000011111111111111111111111101010100011001111100000000000000000000000000000000000000000000000000000000000100000000111111111010100000000000000000000111110101111111111000000000000000000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    28: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011111000010000000101111111111111111100100000000000000010101011000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111100111100111110100000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    29: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101110000001100000111111111111111100110000000000000000000001101100000000000000000000000000000000000000000000000000000000000000000001000111111111000000000000000000000011110011110011111010000000000000000000001111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    30: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000011111111111000111111000111101111111110110000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100100000000000000000001110001111000111110000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    31: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000011111111111111111111111010111001010100100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111110000000000000000000000011100011100011111100000000100000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    32: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000011111111111000000011111111111111011111111111111111011001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110010000000000000000011101001111001011110000000000000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    33: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000001001000000000000000011111111111000000000101011111111110111111101010111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111111000010000000000000001111000111000010111100000000010000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    34: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000111100000010000000000011111111010000000101111111010111111111111110010000011101101111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000011100011110001111100000000000000000000111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    35: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001100000011010000000000000000111111111110000011111111111111111010110101111111010000000111111101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000001110001111000010111000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    36: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001110000001100000000000000000110110111111000001110111111111111110000010001111111100000000010111111111110111010000000000000000000000000000000000000000000000000000000000000000000000000001111110000100000000000000111100011100001111010000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    37: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000110000011111000000000000000111111011110100010101001011111111111000000000010111110100000000000111111111011111101000000000000000000000000000000000000000000000000000100000000000000100000111111000000000000000000010110001111000011101000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    38: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000110000001110000000000000000111111111110000000000000101110001011110000000000001111110000000100001011111111111111111101001000010100100100100000000000000000000010000000000000000000000000001111110000000000000000001110001111100011110100000000000000100111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    39: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001110011000001111000000000000001111111111111000000000000001011100101111010000000000110111000000000000101101010111111111111111111101011011011011101111000100000000000000000000010000000000000000111101100000000000000000011100011101000111000000000000010000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    40: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011100000111110001000000001111111111110000000001000000111100000011100000000000000111111000000000010000010100010110111111111111111111111111111101111011010100000000000000000000000000000000001111101000000000000000101010000110000011110100000100000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    41: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011000000000011000110000011101000010000010111111111111000000000000000011110010001111100000000000001111100000000001000000001010011001010101011011011101101111111111111101101000000000000000000000000000000000011111010000000000000001011000111110001111000000000000000001111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    42: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010100100000111011010100011110000000000011111110111111000000000000000001110000001010110100000000000011110000000000000000000001001000100100000001000000100000101011101111111110100000000000000000000000000000001111101000000000000000011100011101000111100000000000000000111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    43: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000001100110000011111110000100111111011111101000100000001000000111000000011101000000000000001011010000000000000000001111111111011111010000010000000000000010111111111011010000000000000000000000000000111110010000000000000001110010111000011110000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    44: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000001110101100000111111101000001111111111110000000000000000010111100000000011100001000000000101100000000000000000100000111111111111101111000000100000000000000010111111100100000000000000000000000000001111100000000000000000010000111110000111100000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    45: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000100000110100110000111111111111111111111101111000000000000000000001100000000000010000000000000000111110000000000000000000000011011011111111111110000000000000000000010111110111001000000000000000000000000011111100000000000100111100011111010110100000000000001011111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    46: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000000000000011100000000011110111000111111101111101111111111110000000000000000000101110000000001000000010000000000010111111010000000000100000000001011011111111111111100000000000000000001111101100000000000000000000000001011110100000000000000001100001011000011110000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    47: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110110000000000101100001000001101011111111011111111111111101110110000000000000000000011100000000000000000001100000000001101111111110100100000000000000000000001011011111111010000000000000000010111111010001000000000010000000000111111000000000000000110000111100011110100000100000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    48: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000100000111000000000111111011111111111111111101111111101000000000000000000000110000000000000000010111000000000011111111111111010101001000000000000000000111110111111100000000000000000010111101000000000000000000000000011111000000000000001011000011110000111000000000000010111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    49: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000011100000000000111110111111110111111111111110111000000000000000000000100000000000000000010011110000000000000010111111111111101010100000000000000000010111111111000000000000000000011111100000100000000000000000000111101000000000000011100001111000011110000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    50: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000100001110100000010011111111111111111111111111111010000000000000000000000000000000000000000000010111000000000000000000000101011111111111010000000000000000000111111111000000000000000000111111000000000000000000000000111110100000000000001110000111100001110000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    51: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000011000000000000111111111111111111111110101010001010101000000000000000000000000000000000001111110000000000000000000000000101111101111111010000000000000000111111101000000000000000001111110000000000000000000000001111000000010000000110000011100010111000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    52: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110000000000000111000000000000010111111110110111111000001011111111111010000000000010000000000000000000001110100000000000000000000000000000011111111111100000000000000001011111010000000000000000001110100000000000000000000000111110000000000000011100001111000111110000000000101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    53: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101000000100000001101010101001011111111111111101101010101101111111111011010000000000000000001000000000000111110001000000000000000000000000000001011011111110000000000000000111111100000000000000001011111000000000000000000000011111100000000000010101000111000001110000000000110111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    54: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000101111111111101111111111000100101111110100000001011111111101000001001010000010100001000011111000000000000000000000000000000000001011111011100000000000010011111111000000000000000101101100000000000000010000001110100000000000001100010111100001111000000000011101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    55: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000100000010010111111111111111100000000011101000010011111111111111011111110110111111110010100000000111110000000000001000100000000000000000000011111111100000000000000011111110000000000000010111100001000000100000000000011010000000000000111000011110000111010000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    56: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111110000100000001101011110110110101000000110110000001110110111011111111101111111011111011111111101000001111010000000000000000000000000000000000000101111111000000000000000101111100000000000000010111100000100000000000000111111000000000000011000000111000011100000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    57: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101111101011110111111111111111111111010000000000111000001111111111111101111111111011011101111111111101111101000011110101010000000000001000000000000000000001001111110000000000000010101101000100000000001111110000000000000000000000111100000000000001110000111100001111000000001110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    58: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111101111111111111111101000000000101110100110101000111111111111111101000100100101011111111111111110101111101011111101000000000000000000000000000100111111000000000000000111111000000000000000010111000000000000000000010011110000000000001010010011100001101000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    59: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111010010000000000111100000011000111111111010111110000000010110010000010111101111011111011111111110110111001000000010000000000000000001111101000000000000010111110000000000000001111100000000000000000000101110000000000000111000001100000111100000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    60: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011111101110111111111110100100000000001001111100000000011010101000010110100000010011111101101000000111111111101111111111111111111110101000000000000000000000001011110000000000000001011110100000000000000011111000000000000000000010111010000000001001000001110000010110000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    61: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111010101000010000000000000000110110000001001111110100010011110000011011101111111101010000000011111111111111101011111111111111110000010000000000001001111111010000001000000000111101000000000000001111100000000000000000000111000000000000011100000111000011011000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    62: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101001000010101010000000001011100000000111111000000011011010101111111110111111111110000001001111111111111101011111111111111111010000000000000000111101111100100000000000000111110001000000000000111110000000000000000000011110000000000001110000011000001110100000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    63: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111000000101110000000111111000000000101110100011111111110011111111010000100000011111111111111111011111111111111111010000000000000011111111110000000000000000001111100000000000000011111000001000000000000011110000000000000110000101100000011000000011011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    64: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111110000010110000001001111100000000001111100000111111111011101101000000000000000000001011011111011111101110101111111101010000000000011111110111000000000000000000111110000000000000000111110000000000000000000111100000000010011000001110000011110000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    65: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110101111111000001010000000111101000000000101110100011111111111110110000000000000000000000000101111111111111110110111111111111011000000000111111111111100000000010000000001111000100000000000011101000000000000000000011100000000000011100000110000000110000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    66: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010111101000111000000001111100000000010111100000011110111111100000000000000000000000000000000111111111111111100000111111111111110000000011111111111111000000000000000000111100000000000000001111000000000000000000011100100000000001100000111000001011000000111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    67: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000111111110001101000001111100000000000101110010001111011111110000000000000000000000000000000000101001111111111110000010111111111111100000001111111111111100000000000000000011110000000000000001111110000000000000000001110000000000001110000011100000111100001011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    68: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000110000000111010000000010111111000011111111111110000000000001000000000000000000000110001100111111111100000111111111110110100011110111101111111000000000000000001111100000000000000011011000000000000000000111000000000000111000001110000001100000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    69: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100101001001011111000000000011111000001011111011111111000000010010000000000000010000000010101100011111110100000001111111111111100001111111110011111110000000000000000111110100000000000011111110000000000000000111100000000000011100000111000000110000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    70: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110111000000000001111010000000001011110000111111100001011000000000000111000000000000000000001010011100001111111010000001011101111111111000111101110101111111000001000100000011010000000010000001101000000000000000000011100000000000001100010101000000111000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    71: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110100000000001101100000001011111000011011110010000011000000000000011000000000000000000100100010100000011111100000000111110011111111101111111110001111111110000000000000001111000001000000000011111000000001001000001110000000000001100000111000000011000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    72: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001011111000001000011110100101111101000000101100000000000001101000000000000000001010011000000101111111010000001111000011111110101111111000001111101100000000000000111101000000000000011110100000000000000001011000100000000110000001100000001100001110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    73: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111011111010000000000111110000000011111100000111110100000000101000000000000101000000000000000000001010011100000000111111000000000111010011011111111111111000000111110100000000000000011100000000000000001111100100000000000000111000000000000011000001110100000110000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    74: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011011000000000101101000111111110000000001100001000000000001100000100000000000001010110000000000011111100000000111100001111111111111111100000011111110000000000000001111000000000000000111110000000000000000101100000000000001000001010000000110010111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    75: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101000010000101110100000001111010001011110100000000010100000000001000001000100000000000000001100011100000000001111110000000001110000111111111011111000000001111111100000000000000110000000000000000011110000000000000000111000000000000000000000111000000011001011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    76: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001111110110000000000011110000000011111000011111101000000000001001000000000000000100000000000000000001110111000000000000011011000000001111000001110111110111110000000011111101000000000000111100000000000000000111100000000000000001110000000000000010001010100000001100011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    77: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010111111111000000000001111110000001010100000011111100000001000010000000000000000001100000000000100000001010011100000000000011011100000000111100000111111111111110010000000111110100000000000011110010000000000010111110000000000000001111000000000000000000011100000000010011111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    78: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111110000000000001111000000001111000001101110000000101100000000000000000000000100000000010100000001101111000100000000001100110000000011100000111111111111110000000000111111101000000000001110000000000000000011110000000000000000101000000000000000000001110000001010001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    79: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111011000000000000011101000010111110001011111000001001010000000000000000011100111000000000011100000000110011100000010000000101010000000101110000001111111111111000000010001111100000000000000011000000100000000011110100000000000001011000000000000000000000110000000001011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    80: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111111111101000010000001011110000000011000000111111100000001111000000000000000000111101100000000001100000001011011100000000000000010101100000011111000000011101111111100000000000111111000000000000110100000000000000000111000000000000000111100000000000000000000101000000001000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    81: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010011011111111110000000000000011100000001101000000111110000000011100000000000000000000011110000000000001100000001001011110000000000000010000100000000111100001011111011111110000000000011111101000000000011010000000000000000111110000000000000001110000000000000000000011000000000100111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    82: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111011111000000000000001111010000111100000011111010000001111000000000000000000000000000000001000001100000000110001100000000000000001010000000000011100000001111111101101000000000001111101000000000001101000000000000000111110000000000000001100001000000000000000001100000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    83: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000011111111111111111101000000000000111000001011000001111111000000110100100000000000000000000000000000000000001100000000011000110000000001010000000000000000001000000000111111111110000000000000111111000000000001110000000000000000001110100000000000101010000000000000000000010100000000000011011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    84: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001110111111110101111100000000000001100000101111000000011101001000011110000001000000000000000000000000000000000110000000001101011000000101111110000010000000000110000000001101111111100000000000001111110000000000011000000000000000001111000000000000000111000000000000000000000110000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    85: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101101111111111010011111000000000000001110000011100000111111110000001110000000000000000000000000000000000000000000011000000000100011000000011111111100000000000000000000000101111111111010000000000010111101000000000011010000000000000000111110000000000001011000000000000000000000011000000010011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    86: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111111010000011111000000000010011100001011000000011111110000101110000000000000000000000000000000000000000000101000000000100011100000011100111100000000000000000000000000111111111110000000000000111111000000000011000000000000000000011010000000000000111000000000000000000000001000000000001111010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    87: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111010000001011111000001000000011010001110000101111111000000111000000000000000000000000000000000000000000000011000000000110001100000011010001110000000000000000000000000001111111111010000000000011111100000000001110000000000000000101110000000000000010100000000000000000001011000000000000011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    88: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111100100000000111110100000010000111000101110010011111110100001110100000000000000000000000000000000000000000000001100000000010001110000011110011110010000000000000000000000010110111111100000000000000111111000000001010000000000000000011111100000000000001010000000000000000000000110000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    89: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000100000000000111110000000000000111000110100000011111110000101110000000000000000000000000000000000100000000000000110000000011001110000000111111110000000000000000000000000000011111111111100000000010111101010000001011000000000000000000110100000000000011100100000000000000000000001000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    90: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000111111000000000000110001011000001111111000000111110000000000001000000000000000000000000000000000000101000100001001111000010110110100000000000000000000000000000001011111101010000000000011111000000000010100000000000000000111100000000000000110000000000000000000001000000000000000111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    91: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011110000000000011100011110000010111110100101111000000100000000000000000000000000000000100000000000110000000011010110100000011010000000000000000000000000000000000111111111111001000000010111100000000011000000000100000001011110010000000001100000000010000000000000101000000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    92: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000001101001100001011111010000001111100000000010100000000000000000000000000011010000000011000000000100111000000000001000000000000000000000000000100000000101111111110000000001111111000000000000001000000000000101101000000000000111000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    93: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000010100111100000111111100000111111100000000010100000000000000000010000000111010000000001000000001010111100000000000000000000000000000000000000000000000010101111111100000000101111000000001100000000000000000001110000000000000011100000000000000000000000000000000000000011111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    94: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000101111110000000000111001110000001111100000000101110100000001010100000000000000000000000001011101000000011000000000110011110000000000000000000000000000000000000000000000000010011111000000000111111000000000100000000000000000001111000100000000001000000000010000000000000000000000000100011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    95: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111010000000000111001110000111110110000011111111000000001010000001000000000001110000001100011000000101000000000010011110100000000001000000000000000000000000000000000000000100101100000000010111100001000010000000000000000001111100000000000011010000001001000000000000001000000101110101011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    96: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000111111100000000001110011101000011111000000001111111100000101100000000000000000000111000010100001110000011010000000011001111000000000000000000000000000000000000000000000000000000000000000000001111110000000100000000000000000000111100000000000000100000001110100000000000000000000111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    97: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010110101100001101111000001011111110100000011000000000000000000000010000000110000011000011000000000001100111110000000000000000000000000000000000000000000000000000000001001000000111111001000010000000000000000000011110000000000001010000001111111000000000000000001111111111010111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    98: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000011011111100000000011010110000010111100000000111110111000001101000000000000000000001110000010010000101100010000000000001100111000000000000000000000000000000000000000000000000000000000000000000010111110101110000100000000000000000011110000000000000100000000111110100000000000001001111111111010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    99: dataREG =  641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011111111101000000011101111000101111100000011110111111000000100000000000000000000001110000001100000011011100000000000001010111110000000000000000000000000000000000000000000000000000000000000000000011111111111010000000000000000000011111000000000000111000000011111000000000000000000111111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    100: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111100001000111111110001011111100100001111111110100001110000000000000000000000101000001010000000110000100001000000110001110101000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000111100010000000010000000111111110000000000000000111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    101: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111101111100000000111111100001111111000000001111110110000001000000000000000000000010110000000110000000001000000000000000010011111000000000000000000000000000000000000000000000000000000000000000000101111111111111001000000000000000001110100000000000001000000001111101000000000000000011111011111101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    102: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000101000000000111111111111100000010111011010001111101000000111111110110000111000000000000000000000000110000000110000000000000000000000000111001111000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000111100000000000001000000011111110000000000000000111111111111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    103: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000010101001111011000000001111111000001111110000000111111111000000010100000000000000000000001110000001010000000000000000000000000010010111100000000000000000000000000000000000000000000000000000000000000000001111101111110100001000000000000000111100000000000000100000001111110100000000000000011111111011111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    104: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011110101111111100000011101111000111101110000000110111101010000011000000000000000000000000111000000111000000000000000000000000011001111010000000000000000000000000000000000000000000000000000000000000000000111111101111111100000000000000000011111000000000000000000010111111000000000000000011111111111111111011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    105: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111011111110011111111100000001110110000111110100010001111011111100000001000000000000000000000000011100000101000000000000000000000000001100111110000000000001000000000000000000000000000000000000000000000000000000011111111111111000000000000000000001100100000000000000000001101111100100000000000001110111000011111111011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    106: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000111111111100001111011110000111111010000001111111110100010110000000000000000000000000001110000100000000000000000000100000010100011111000000100000000000000000000000000000000000000000000000000000000000111111111111101110010000000000000001110001000000000000000001111111100000000000000001111111101011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    107: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000111011111000000011111100001111111000000010111110111001000011000000000000000000000000000010111010000010000000000000000000001100111110000000000000000010000000000100000000000000000000000000000000000000011111111111111110000000010000000001111100000000000000000000111111110000000010000001111111000001011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    108: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001101111111100000110101010001111111000000011111111111100000101001000000000000000000000000101101000000000000000000000000000000110001111100000000000000000000000000000000000000000000000000000000000000000010111111101111111000000000000000000111000000000000000000000111011110000010000000000111111100000110111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    109: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011110111111010001110111000010111110000000011110111011100000001100000000000000000000000000000101000010000000000000000000000000110101110100000000000000000001000000000000000000000000000000000000000000000011111101110111111100000000000000000011100000000000000000000011111111000000000000001011111110000001010111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    110: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011010111111100001110111000011111100000000011111101110100000010100000000000000000000000000000000001011000000000000000000010000110011110000000000000000000000000000000000000000000000000000000000000000000001011111110011111110000000000000000001100000000000000000000111110111100000000000000101111110000000010111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    111: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101111000011111000001110111000111111110000000111010111010000000001111000000000000000000000000000000000101000010000000000000000000110000111000000000000000100000000000000000000000000000000000000000000000000001111111010001111101000000000000000011110000000000000000000011111111000000000010000011111101000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    112: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111100000111111100011010110000111111000000001011111111110000000000111100000000000000000000000000000000110000000001000000000000000001001111010000000001001010100000000000000000000000000000000000000000000000000111111101001111111000000000000000001101010000000000000000001111111110000000000000011111110000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    113: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110100000111111100001100111000011111100000000111101111000000000000001000010000000000000000000000000001110000000000000000000000000110000111100000000000000111010000000000000000000000000000000000000000000000000111111110000111111100001000000000000110000000000000000000001111111011000000000000001111111000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    114: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000110111000111110100001111111000000001011110110100000000000101000000000000000000000000000101111000000000000000000000000000011000111100100000000011001111000000100000000000000000000000000000000000000000111111101000011111100000000000000001110000000000000010000101111111110001000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    115: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000111111000011001110001111101100000001111101111000000010000110000000000000000000000000000010100100000000000000000000000000101000111100000000000001111111100000000000000000000000000000000000000000000000111111110000101111110000000000000000111000000001000000000001110111111000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    116: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000111111100111101100010111110000000001111110110101000000000110100000000100000000000000000000000000000000000000001000000000001000011110000000000011111000111000000000000000000000000000000000000000000000101111010000001111110000000000000000111100000000000000000000111111111100000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    117: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101101011100010000000000000111111100011001100011011111000000000111111011000000000010100000000000000000000000000000000000000000000000000000100100000010100010100000000000001111001101000000000000000000000000000000001000000000000111111111000001011111000000000000000011010000000000000000000111111111110000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    118: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111011010000100000110110100111001100001111100100000001111111101000000001001100000000000000000000000000000000000000000000000000000100000000010000111110000000000000110100111000000000000000000000000000000000000000000000011111010000001111111000000000000000111000000000000000000001111111101110000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    119: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110101000000000111111001101011000011111110000000001111001110000000010001100000000001010000000000000000000000000000000001000000010100000001000011100000000000000011011111100000000000000000000000000000000000000000000011111110000000011111000000000000000011110000000000000000000011111010111000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;        
    120: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000011111100110001100011111110000000001101110101000000011010110000000001100000000000000000000000000000000000000000101000000000000011110000000000000001111000100000000000000000000000000000000000000000000010111111000000011111110000000000000011100000000000000000000101111110010110000001000001011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;        
    121: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111111010111111111101000111111001110001000001111110000000000101110100000001011011000000000001100100000000000000000001000000000000000000000100000000000011111000000000000001110011110000000000000000000000000000000000000000000011111111000000001111010000000000000101110000000000000000000010111110011010000000000000111011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;        
    122: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000101111111100111111001110101000111111001000001000000010000000000110011100001000001110000000000000000010000000000000000000101100100010000000011000000000000000000111011110000000000000000000000000000000000000000000011101101000000010111100000000000000011101000000000000000000111111111001100100000000000011111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;        
    123: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000010111111111011111001110010100011101110000000000000000000000000110001000000000001100000100000000000000000000000000000000000010100000000000011110000000000000000110101101000000000000000000000000000000000000000000001111110000000001111110000000000000010110000000000000000000011101110101111000000000000101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;        
    124: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001111101111111100000000111111111011101110011000011111100000000000000000000000001010011100000000000100000000000000000000000000000000000000101011000000000100101100010000000000000011010010001000000000000000000000000000000000000000000011111000000001111111000000000000001110000000000000000000001111111100110000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;      
    125: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111011110100000000010111111110101110101000011111100000000000000000000000000110001100000000000110000000000000000000000000000000000000100101100000000000011100001000000000000011100010000000000000000000000000000000000000000000000011111100000000111110000000000000011011000000000000000000001111111110111100000000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ; 
    126: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110011111100000000000101111111101100110100011111100000000000000000000100000110001100000000010110000000000000000100000010000000000000010011100000000000111100000000000010000010001010000000000000000000000000000001000100000100000010110100000000111111000000000000001110000000000000000000001111111010011110000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ; 
    127: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110100111110000000000011111111011100011000111111000000000000000000000000000011001100000001000100000000000000001011010000000000000000101110000000000000011000000000000000000001100100000000000000000000000000000000000000000000000001111000000000110111000000000000011111000000000000000000001101111111001110000000000000011111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ; 
    128: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110001001111000000000000011111111100110000011111110111010000000000000000000101000100000000000110000000000001000111101000000000000000010011100000000000111100000000000000000001111110000000000000000000000000000000000000000000000001111010000000011110100000000000000110000000000000000000000111011101010111100000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ; 
    129: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010001100111100000000001011111111100111000001111011011010000000000000000000011100111000000010110000000000000001110100100000000100001011011100000000000011100000000000000000000011100000000000000000000000000000000111000000000000000111100000000111111000000000000001111000000000001000000000011011101100011110000000000001111110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ; 
    130: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111100000110010100000000000011101111100111001011111111111100000000000000000000001100010000000001000000001000000000111101100000000000000010101100000000111110000000010000000000000010000000000000000000000000000000001011110000000000000111100000000011111001000000000001111000000000000000000001111111101110001010000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ; 
    131: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000001000100000000000011111011000101000011111111111100100000000000000000000101011110000111010010000000000000111101100000000000010110111000010010111100000000000000000000000000101000000000000000000000000000001110111000000000000011110000000111111000000000000001111010001000000000000000010011110111001101000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ; 
    132: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000100001011000000000101111111100111000011011111111000000010001010000000000110000101111110000000000000000000111010110000000000010101011100000011111010000000000000000000000000000000000000000000000000000000001110001100001000000001110001000011111100000010001000111000000000000000000000011101010001000011000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ; 
    133: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111100000101000010001000000111111110100011000001001111110100000000000011110000000010000101011010000000000000000000111100010100000000010110101100001111111100000000000000000000000000000000000000000000000000001000000010001110000100000100111000000011111000000000000000111000000000000000000000010101101011100001100000000000011111000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;    
    134: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000010001010000000000011111111000011000000001111110000000000000011110000000001000000000000000000000000000000011101000000000000010110110100001110100000000000000000000000000000000000000000000000000000000000001101000110000000000001110000000011101000000000000001111000000000000000000000011001111101110000110000000001011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;          
    135: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000000001001111000000000111110110000111000000011111100000000000000101111100000000000000101000000000000000000000111100100001010000011010111000010111000000000000000000000000000000000000000000000000000000000000000110001010000000000000011000000101111000000000000000111000000000000000000000001101110100110000010000000000111111100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;          
    136: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000100100100100000000011111111100001000000111101101010000000000010001100000000000000000000000000000000000000011010000001111000001111011000001110000000000000000000000001000000000000000000000000000000000000000001111110000000000000010100000011111100000000000000111100000000000000000000001100011110011001001100100000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;           
    137: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110110000000000000110101000000101111111000111000000011110000100000000000001000110000000000000000000000000000000000000011100001011010000000001011000011101000000000000000000000000000000000100000000000000000000000000000000101000000000000000000000000001011000000000000000110100000000000000000000001110111111011000001110000000001111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;           
    138: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001111100000000000000000100000100111111101000011000001111111011010000000000110101101000000100000000000000000000000000000000001000011110100111110010000011100000000000000000000000000000000000000000000000000010000000100000000010100000000000000000000000011111000000000010001011000000000000000000000000110001101001100101111010000011011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    139: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000111111100000000000000000010100000111110110000010100000111111001000000000000011010100000000000000000000000000000000000000010000001111110000000101001000011110000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000001111100000000000000111100000000000000000000000110011011010110011111110100001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    140: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000001000000010000000110111111000001000001111110001100000000000001101100000000000000000000000000000000000000000000000111111000001010000000111100010000000000000000000000000000000000000000000000000000010111100000000000000000000000000000000000111100000000000001111000000000000000000000000011000110100110111111111010001111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    141: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000011111100000000000000000000000000111111110000101000001111110101001000000000000110100000000000000000000000000000000000000000000011010110000000001000000111110000000000000000000000000000000000000000000000000000000000111110100000000000000000000000000000001011110100000000000111100000000000000000000000011000011010011011111111111000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    142: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000111111110000011000001111110101001000000000000000000000000000000000000000000000000000000000010111100111000000000000001111100000100000000000000000000000000000000000000000000000000000011111010000000000000000000010000000000111010000000000000111000000000000000000000000011100101100011011111111111111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    143: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010111111000000000000000000000000000111111110000010000011111010011001100000000000000000000000000000000000000000000000000000001011110000110000000000000110111000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000100011110000000000001010000000000000000000000100110000011000001101101111111100111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    144: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000111111101000001100000111100110001100000001000000001000000000000000000000000000000100000000101100010111000000000000011101100000000000000000000000000000000000000000000000000000000000011111101000000000000000000000000000000011110000000000000111000000000000000000000000001110000110001010111111111111111111000111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    145: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110110000000000000000000000000001011111110000101000011111100111000110000000100000000000000000000000000000000000000000000011111000000011100000000001111110100000000000000000000000000000000000000000000000000000000000001111111010000010000000000000000000000101111000000000001111000010000000000000000000011010001000000101011111111111101111100001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    146: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111000010000000000000000000000000110111100000011000011111100100010100000010100000000000000100010010101001000000000010011111101000000011100000001111110111000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000011111100000000000111000000000000000000000000001101000110000101011101111111111110100001111110101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    147: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000111111100000000000000000000000000001111111010000001000011110101110001010010011100000000010000011101111111111100100000000011111000000000001111111110110110010000000000000000000000000000000000000000000000000000000000000001111111100100000000000000000000000000001111000000000001110000000000000000000000000000110010001000010001111111111111011000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;         
    148: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000100000000000000111111110000110000011111001010000111000001010000000000011111111101111110110000000101111110000000000000111111111111000110000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000001111110000000001011000000010000000000000000000111001000000001110111111101111111110000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ; 
    149: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110100000000000000000000100010001111101010000011000101111001100000011000011101000000000011110010110101010000000111111101000000000000000000101110101000110000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000111110000000001110000000000000000000000000000001011100000000011111111111111111000100000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    150: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000001111111010000011000111111001100000001111010000000000011110001000000000000000000111101100100000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000100101000000000000000000000000000000010110110000000000110000000000000000000000000001111011100000000001111111111111111100000000111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    151: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111110000000000000000000000000000011111111000000010000011110010110000011110111000000001011101000000000001010000010110100000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000001111111000000001110000000000000000000000000000010101110000000010111101111111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    152: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111000000000000000000000000000000101101111110000011000011111001000000000001000000000101111000100100100110111000000011100000000000100010000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000011110100000000111000000000000000000000000000011101110100000001101111110111111100000000000111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    153: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000011110111000000001001011111011100000000000000000000101100000011111111011111100000011100000000000010010000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000111110100000010100000000000000000000000000000000100111000000000111111010101111110000000000011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    154: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000111111111100001010000110110011000000000000000010011110100000111111111111110000000101100000000000000011100010000010111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000011111100000001110000000000000000000000000000010110111100000000111111101111101110000000000001111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    155: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000111111111100000111000111110001100000000000000000101110000000110100101000111100000011100000000000000000111000010101000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000010000000000000000000000000000001010111000000000101111100011111101000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    156: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000011011111111000000000000111111011000000000000000001111000000010111000000000111000000011100000000000000010101001011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000100000000000000000000000000000001010111110000000011111110001111110000000000000101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    157: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010000000000000000000000000000011111111111100000111000111100001100000000000000101111000000001101000000000011100000011100000000000000000001001101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000010000000000000000000000100000001010011101000000111111010000111110000000000000011101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    158: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011000000000000000000010000000000111111110110000000101000111110010100000000000001110100000000111100000000000110100000011100010000001000000000001110101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111101000000000000000100000000000000010000000010111100100000011111100000011110010010000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    159: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000001000100001011111111011111000000010001111101010000000100000010111000000000011010000000000011000000011101000000000000000000111100010000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000001011110000000000000000000000000000000011000000001001110000000011011110000000101000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    160: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001111111000001000000000000011011110111110111111111010000111010111100001100000000000011110000000001111000000000000111100000011100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000010100000100011111000000001111110000010000000000000000000010111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    161: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111110000000000010000000001110011111111111001111000000010001111110010000000000000011010000000001110000000000000011010000011000000000000000000000001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000010100000000001111100000001111110000000000000000000000000001101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    162: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010000000000000000000000000000011111010001101000000110011111100010000000000001111000000001111010000000000000011100010111000001010000000000000011110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000001100000000001111000000101110110000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    163: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111101101000000000000000000000000000111111110111110000000110010111100001100000010001011000000101111000000000000000001111011111000001100000000000000011101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000110000000001111110000001111101000000000000000000000000000011101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    164: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111100000000000000000000000000101111111000001111000000011011111110010000000101001111000000011101000000000000000000111111100000000010000000111000000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111000010000000000000000000000000110000000000111111000001111110000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    165: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000111101110100011110010000101011111100000000000010000111010001111100001000000000000000011101110000001100000000101000001100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000011000100010111111110000111111000000000000000000000000000001111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    166: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000100000011111111111010000111110000000111011111010000000000011001011000000111010000000000000000000010100000010011010000000110000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000111000000000110110111111111100001000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    167: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000001011111111110100000101110000001010110111000000000000110100110000000111000000000010000000000001010000000011000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000010000000011000000000111111110111111111000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    168: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000001111111111110000000111111000000111011111000000000000011000111000000011000000000000000000010000000000000011000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100010000000000000001010111010000000000000000000000000000001110000000011111111011111111000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    169: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101111100000000000000000000110111010000000010111111000000101011111000010001010011000111010010011100000000000000000000000000000001101000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011001000000000000000111111110100000000000000000000000000001010000000110111111111101110000000000000000000000001000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    170: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111110110000000000000000000010101000000000001111111000000111011111000000000101011001111100000111100000000000000000000000000101010100000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111000000000000000011111110000000000100000000000000000001110000000010111111111111111000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    171: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101100100000000000000000000000010000000011111011100000010101111000000000111011101111000000011100000000000000000000000000111111100000000000111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111101111100000000000000011111111010000000000000000000000000001010000000011101111111111110000000000000000000000000000000000001111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    172: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101110000000000000100000000000000000000101111111000000011011110100000000011111010111110000001110010000110000000000000001101010000000000000001101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011111000000000000000101111111100000000000000000000000000000111000000010111111111111111000010000000000000000000010000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    173: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000110000000000000010000000000000000000011111111110000011001111000000001011111111111010000001110000000110100000000000010100000000001000000011110101101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100001111100000000000000001011111110000000000000000000000000000011000000010111110110111111000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    174: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111000110000000000000000000000000000000001101111111100000011001111100000000111111111111100000100110000001010000000000100011100000100000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111010001111100100000000000001111111110001000000000000000000000000111010000010111111111111111100000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    175: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010001111000000000000000000000000000000000111111011100000101011111100000000111111011111101000001111000000110000000000011001000000000000000000000001001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000111111110000000000000011110111011000000000000000000000000000101000000011011111111111111000000000000010000000000000000010000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    176: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000111000000000000000000000000010000001111101101111000011100111110000000010111111011100000000111000000110000000000110001110000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110000110000110000000000000000111111111000000000000000000000000000011100000000101111110101111100000000000000000000000000000000000000101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    177: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000111100000000000000000000000000100001111110001111000001000111010100000111111111111100000000011010000011000100000111001100000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111010000110100000000000000111011111100000000000000000000000000001100000011010111110111101100000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    178: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000110100000000000000000000000000000111111100101111000011100111110000000111111111110100000000111000000010000000000100001110000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000011101000000000001111101011110000000000000000000000000010100000001111111111001111101000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    179: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111100000011000000000000000000000000000011111111100011111100001010111100000000011111111111000000000011000000111000000001110001100000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001110000000000000111111101101000000000000000000000000001110000001001111110001110111100000000000000000000000000000000010010111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    180: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000110110000000000000000100000000001110111000001110100001100011111000000111111111101000100000011100000101000000001110000110000000000000000000000010100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000111010000000000011111010111000010000000000000000000011110000011111011111000010011001000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    181: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000010010000000000000000000000000111111010000001111110001100011111100000011101111110000001000011110000111100000000110000111000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001110000000011100000000000111111101011100000000000000000000000001010000001011110110000000001100000000000000000000000000000100010110111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    182: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000101000000000000000000000000001101111100000011111100001100011111010001011111111010001100100011000000011000000001100000010000000000000000000000011000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010101000110000000011101000000000011111110111100000000000000000000000001110000001001111110000000001110000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    183: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111000010100000000000000000000000000111111010000011111110001110011111100000111111111100001111000011100000011100000011100000111000000000000000000000101001010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000011000000001110000000000111111110001110000000000010000000000000110000000010111111000000001101000000000000000000000001011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    184: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000001000000000000000000000000000111100000000001111010000110001111100000001101111000001111111111000000011000000000111001010000100000000100000000110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011100001111111000000000011111111100111100000100000000000000001011000000001111110000000000111000000000000000000000000111011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    185: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111010000100000000000000000000000000100000000000001111111000110000111110000111110111100000111101111100001011101000001100000111000000000000000000000111000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110110101111000000000001111111110111010000000000000000000000110000000000111110000000000111010000000000000000000010111111111010111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    186: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000100000000000000000000000010000010000000000111111100000110000111110000011111111000111101010100000001100000000000111000111000000000000010000000100000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101011111100111000000000111111110100011100000000000000000000000111000000011011110000000000111000000000000000000000011111111011011011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    187: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000010011111111001011001011110000111111111100001110000010000110110000000000011101010000000100001100100001110000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110100000110000000000011011111110011111000000000000000000000110000000001111110000000000101110000000000000000000011111101000000101101110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    188: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000111111110000111000111111100011111111000001110000000000111000000000000000111110000000000010111000000111000000110000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001111000000011100100000001111111110000111000000000000000000000011000000000111111000000000111010000000000000001000111111010100000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    189: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000010000000000000000000000000000001000001010111111000111000101111000011111101000011110000000001101000000001000100101000000000000011101110000111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000011100000000011111101111000011110000000000000000001011000000001111010000000000111111001000000000000000110111100001011100000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    190: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000001110111100001011100011111000011111101000011010000000010100000000101110000001000000000000010101000100101100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000110000000000101111100111000101110000010000000000000011100000000111110000000000111110100000000000000000111110000001101110010001011111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    191: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000100000000000000000000000000000011011110111000111000011011100010110000000011100000000011100000000011111100000000000000000111011000000111011110000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001100000000011100000000011111100111000011111100000000000000000111000000011111100010000000111111000000000000000010111111000010110111000000101001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    192: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111101000000000000000000000000000000000000000101001111110000111100001111110011111000000110100000000001000000001011001100000000000000000001101100000001110101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000011100000000010111010011110000111010000000000000000001000000000111110000000000101111100000000000000001111111100001010001100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    193: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110100000000000000000000000000100000000000111001111110000111100001111110001110000000011100000000011010000000010001110000000000000000001110000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001010101100000000011111100011100000111110000000000000000011100000010111110000000000111111111000000000000000111111100001011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    194: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000000000000000000000000000000000111010011111110000111100001110110011111000001110001001000011000000000011000101000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001100001111110100000000011111100010110000011111000000000000000011000000001110100000000000011111110010000000000000010111110000010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    195: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000101000000101100011111010000111110000111110001100000001111000110100001110000001010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110111111000100000101111000011100000011111110000000000000101100000011111100000000000011111111000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    196: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110100101010000000000000000010110111111010001111111100000111110000111111011110001000110001011100001100000000011111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111010100111100000000011111110001111000001111110100000000000011000000000111110000000000010111111100000000000000000111111000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    197: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111110000001101001000000000000000011100101000000111111100010111101000110110000100101011101001011100000111000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111010000011000000000011110100000101000000111111110010000000001100000011111100000000000011101111101000000000000100011111110000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    198: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000111111000000000000000000000010000000111111111100001111100000111111000000100101100011001110000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000110000001011000000000011111000001110000001111111010000001000101000000011101100000000000001111111101000000000000000001111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    199: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101000010010100000001000000000000000000101011011111010001111110000111111000010101111000101000100000101000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000111000000110000000000011111100000111000000011101111000000000011100000101111100000000000011111111000100001000000000010111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    200: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000101101000000000000000000000000010011110110111000101111110000011101100001110110100011100111000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000011101011110000000000011111000000111100000011111111111000000001000000011111010000000000000111111110010000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    201: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000010111000000000000000000000000011011000111111000010111110000011110100001111110000101000101111110000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111011110000000000011111110000010100000001111111110000000011100000111111100000000000001101101011001000000000000000011111110000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    202: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000011010100000000000010000010111011101000111110000011111110000101111000001111000000011000010111010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101101000010000100101110000000111100000101111111111000000010100000111111100100000000001111111010101000000000000000010111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    203: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001110110000000001010000000000000000000101010101000001111110001111111100000011111100101110100000101000011011000000000000000001000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000000000000111111100000011000000011111011110000000011000001111111010000000000000111110111000100000000000000001111110000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    204: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101000000000000000000000000000000000101000000001111010000011110100000111111100111100000000011000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000011110000000111110111000001000100001011111000000000000001111111001110010000000000000010111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    205: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000101111110001101111110000011101111111110000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000010000000000000000000000000000000000000000000000000000000000000000000000000000111111000000001010000001111111111000000011000001111111100000000000000111011001101001000000000000000011110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    206: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001111111000001000000000010000000000000000000000000000011111000000110111000000011111111010110000000011000000000100000100000000000000000000000000010000000000000000010000000000000000000000000000000001010001000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000011100000000111110111000000101100011111111000000000000000111111000110100100000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    207: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000111111000011001111100000101111101001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000010000000000000000000000000000000000000000000000000000000100000000001111101001000001110000010111111111000000010000011111111100000000000000011101000110000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    208: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111000000000000000000000000000000000000001000000111110100010100111100000011111010000110111101010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010101000100000000000000000000000000000000000000000000000000000000000000000000000000010111111000000001110000001111111111000000011000111010110100000000000000111111100001000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    209: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111100000000000000000000000000000000000000000000010111111001010000011000000011111000000111111111011010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010101010010000000001000000000000000000000000000000000000000000000000000001110000001111110000000001110000000011111111000000101000011111110100000000000000011111000000000000000000000000000010111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    210: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111010001000000000000000000000000000000000000000011101111000110001111000000011111000000011011111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001001000000000000000000000000000000000000000000000000000000000000000000001011000001101111011110000110000000001111111000000011001111111111010000000000000111111000000000000000000000000000111011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    211: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000100000000000000000000000000000001011111111110100000011000001011100000000011110111111111111111111001000000000000000000000000000000000000000000000000000000000000000000000000000000000110010101010000000000000000000000000000000000000000000000000000000000000000000111100011111101111111001110000000001011111000000100000111111111100000000000000011101100000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    212: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100111111111000100000000000000000000000000000000000000000111111111011100100010000000111111100000011010101111111111111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000001001000100000000000000000000000000000000000000000000000000000000000000000000001101011111110111111000111000000001111101000000011001111111111000000000000000001111000000000000000000000001000011111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    213: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101111100010011010000000000000000000000100000000000111111111111111000000011000000011110000000011100110110111111111111111101111010000000000000000000000000000000000000000000000000000000000000000000000000001011001000000000000000000000000000000000000000000000000000000000000000000000000111011111110111111100110000000001110111000000100001111111111100100000000000011111100000000000000000000000100111111111010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    214: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101001011111000010000000000000000000000100000100111011110111110100001010000000111111000000111011010110111111010111111111111011001000000000000000000000000000000000000000000000000000000000000000000000010011001100001000000000000000000000000000000000000000000000000000000000000000000101111111011111110001111000000001111111100000110101111111111000000000000000011111000000000000000000000000001011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    215: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110111111100011010000000000010000010111111011111111111111110000111100100000111100000010111001001001101111010101111111111111110000000000000000000000000000000000000000000000000000000000000000000001001001010101100000000000000100000000000000000000000000000000000000000000000000010011111111111011110000010000000000110110000010000011111111111100000000000010011111100010000000000000000000001111111111111000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    216: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000111111111111111111000101100000000000000000011111111111111111111111100000010110000001111111000001111011101010111011000000010101111111011110100000000000000000000000000000000000000000000000000000000000000001000111011000011000000000000000000000000000000000000000000000000000000001000000000001111111011111111000111000000001011111000000110111110111111000000000000000001111100000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    217: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011101011111111000111000000000000000000011101111111101000011111110000111110000000111110000001000010011001111111000000000000010111111111111000000000000000000000000000000000000000000000000000000000000001010101111101100000000000000000000000000000000000000000000000000001000000000000000000110111111110110000101001000000111111000010000011111101111100000000000000010111100000000000000000000000010111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    218: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000111110000111000000000000000010001110101000000001011111000011111000000001111110000001100101000101111100100000000000010111111111011101000000000000000000000000100000000000000000000000000000010000011111111110100000000000000000000000000000000000000000000000000000000000000000000000111111111111110000110000000000011111000001001111111110111100000000000000011111100000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    219: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110010000000101101011110000000000000000000000000000000000100111111000000111100000010111110100010000100110011111110000000000000000000011011111110100000000000000000000000000000000000000000000000000000000000101110111010000000000000000000000000000000000000000000000000000000000000000000000000111111111111010000011000000000010111000001000111111011111010000000000000011101000000000000000000000000111011010100001110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    220: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010111000000001111110001111100001000000000000000000000000000001111110100001111101000011111110000011000010110111111110000000000000000000100111111111011101000100000000000000000000000000000000000000000000000000011111111101000000000000000000000000000000000000000000000000000000000000000000000001111111101111100000110000000000011001000000101111111100111100000000000000001111100000000000000000000001011110100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    221: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000001111000111110000000000000000000000000010000000000111111000001110100000011101110000001000000000011111110000000000100000000000000101111110100000000000000000000000000000000000000000000000000000000001011111100000100000000000000000000000000000000000000000000000000000000000000000000111111111111110000011000000000011111000010010101111000110110000000000000001111100000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    222: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110100000000011111100111110000000000000000000000000000000000011111100010011111000000011111110000111000001001010111101000000000000000000000000111111111111100000000000000000000000000000000000000000000000000001011101110100000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000110000000000011011000000011111111001111010000000000000001111100000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    223: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000001011111000111110010000000000000000000000000000000011011110000011111000000111111111000001000000000110111100000000000000000000000000000111111111110000000010000000000000000000000000000000000000000000001111010000000000000000000000000000000000000000000000000000000000000000000000010101111111111111100000010000000000001110000101011111110000111100000000000000001111010000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    224: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111000000000111110001111010000000000000000000000000000000000011111100000001111100001111111110000010000111001111111110000000000000000000000000000000111111111110100000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000011110111011110100000101000000000000111000000011111101001111100000000000000001111000000000000000000000101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    225: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000010111010001111110000000000000000000000000000010000111101100000011110100001111111110000011000111100100111110000000000000000000000000000000001111111111000000000000010000000000000000000000000000000000000111101000000000000000000000000000000000000000000000000000000000000000000000000111111111101111100000010000000000000110100110111111100000111110000000000000001111100000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    226: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000001111100111110000000000000000000000010000000000000111110000001011111000101111110111000010000111111110111010000000000000000000000000000000100111111111110000000000000000100000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111010000100000000010000110001000111111110001111110000000000000001111000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    227: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011111000010111100000000000000000000000000000000001111111000000111111000111111111110000101000111111101111100000000000000000000000000000000000001111111111010000000000010000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000010010000000000110000101111111000001111010000000000000011111100000000001000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    228: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100011110000010110000000000000000000000000000000000101111110000011111111010111111111111000011000101111010111110000000000000000000000000000000000000101111111101000000000000000000000000000000000000000000001111110100000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000110010011110111000001011101000000000000000111000000000000010000000011111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                                                                                                                                                                                                                                        
    229: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000111010000000000000000000000000000000000000000000011111010000001111111011011110111111000001000010111100111110010000000000000000000000000000000000000101111111101000000000000000000000000000000000100000100111110000000000000000000000000000000000000000000000000000000000000000000000001010110101111111100000000000000000000110000011111111000001111111000000000000001111100000000000001000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                                                                                                                                                                                                                                        
    230: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000001000000000000000000000000000000000001101111100000101111111011111111111110100010000011111010111110000000000000000000000000000000000000010111111111101000000000000000000000000000000000000000001110110000000000000000000000000000000000000000000000000000000000000000000000000011111011011111111000000000000000000010000011111110000011111110100000000000001111000000000000101000000111111000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                                                                                                                                                                                  
    231: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110100010000000000000000000000000000000000000010111110000100111111011111110101110111000011000000111001111110000000000000000000000000000000000000000001111110110100000000000010000000000000000000000000000111110100000000000000000000000000000000000000000000000000000000000000000000000000110011111111111100000000000000000100000111111110000001111110000000000000010111100000000000011110000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                                                                                   
    232: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111010000000000000000000000000000000000001001101111011000001111011111111111010111101000001000000101110111111000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000011101111111111100000000000000000000000111111100000011111111100000000000001111000000000000001101000011111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    233: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101000000001000000000000000000000000000101111111100000101111111111111111101111111000000100000110010111111100000000000000000000000000000000000000000001111111101100000000000000000100000000000000000000011110000100000000000000000000000000000000000000000000000000000001000000000000000011101101111111110000000000000000000001011011110100010111111100000000000001111100000000000000111100101111100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    234: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000001000000000000000000101111111111110000000111111111111111111110111111000010000000111001111111000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000001011100101011111110111111100000000000000000000000111110000000111110111100000000000001101000000000000000101100111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    235: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111100000000000000000000000010000010111111101000000001111111111111010111111111110100001000000111000111111100010000000000000000000000000000000000000000010111111111010000000000000000000000000000000000101101000000000000000000000000000000000000000000000000000000000000000001011111011111111101111011110000000000000000000000011111000001011111110100000000000001111000000000000000011111110111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    236: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111000000000000100000000000000111111010010000000011101101111111101111111111111000000010000011110111111110000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000111110000000000000000000000000000000000000010000000000000000000000000101110111111111111010101111100000000000000000000000111110000000111111111000000000000010111100000000000000000110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    237: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010000000011111100000000000000000000000000001001000000000001111111101010101000011110111111000000000000011100110111110000000000000000000000000000000000000000000000011111011111100001000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000010111111111111101111000010111110000000000000000000000111110000001111111110100000000000001101000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    238: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111000000000001111010000000000000000000000000000000000000000011111111001011110001011111011111100000001001011110111111110000000000000000000000000000000000000000000000001111111110100000000000000000000000000000000111010000000000000000000000000000000000000000000000000000010000000011111111111101111110000001111110000000000000000000001111100000011011111110000000000000011111000000000000000000001111101110000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    239: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110100000000000111100000000000000000000000000000000000000010110111000000000110000111101111111000000000000011000111110111000000000000000000000000000000000000000000000000101111111110000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000001101111110111111111111000000111100000000000010000000010111010000001111111000000000000000001111000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    240: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000001110000000000000000000000000000000000000001111101100000001111000011111111111100000000000001110110111111100000000010000000000000000000000000000000000000011111111111100000000000000000000000000000111100000000000000000000000000000000000000000000000000000000001011111111011111111111100000000011111000000000000000100011101100000011110111110000000000000001111000000000000001000000001111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    241: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000011111000000000000000000000000000000000000111111100000000001101000011111111111110000010100011100111011111101001000001000000000000000000000000000000000000001111111111110000000000000000000000000000111110000000010000000000000000000000000000000000000000000000001111111111101001111111110000000111110000100000000000000011110000000111111101000010000000000001110100000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    242: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000001111000000000000000000000000000000000010111110000000000001110001011100111111000000000100001100111011111110000000000000000000000000000000000000000000000110111111111111000000000000000000000000000111100000000000000000000000000000000000000000000010000000000101111111001111100111101110000010011111000000000000000001111111000000111111110000000000000000010111000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    243: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110000000000010011111000000000000000000000000000010000101110000000000000001110000011110001111110000000000001000010011111110000000000000000000000000000000000000000000000111111111101111100000000000000000000000000111100000000000000000000000000000000000000000000000001000011111111100000111111111111100000000111110000000000000000111111110000001111111100000000000000000011110000000000000000000010000000111111010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    244: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000111110000000000000000000000000000000011001000000001000011111000001110111111100000000000001100011000111111100000000000000000000000000000000000000000001011111111111111111000000000000000000000000011010000000000000000000000000000000000000000010000000001111111111011000011111111011100000000011111000000000000000001111111000000111111110000000000000000001111000000000000000000000000000011111100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    245: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000010000100000001111000011110111111110000000000000101011001011111110000000000000000000000000000000000000000001111111011111011111100010000000100000000000111110000000000000000000000000000000000000000000000000011111111101000100001111111101110000001011111100000000000000111111110010011111111000000000000000000010110000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    246: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000011000011101000001111011111110000000010010100011000111111110100000000000000000000000000000000000001011111111111111111011110000000000000000000000111000100000000000000000000000000000000000000000000111111011110000000000111111111111000000000111111010001000010000011110110000011101110000000000000000000011111000000000000000000000000000000111111000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    247: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000111000001110000011110110111101000000000001010011000011111011000000000000000000000000000000000100001111110111111111111111010000000000000000000001011110000000000000000100000000000100000000000000111011111111001000000000001110111111101000000011111100000000011100001111100000111111101000000000000000000011100000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    248: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011100000000000000000000000000000000000000000000011000001111100001110001111110000000000000100001100000111111110000000001000001000000000001000000101111111111111111011111111100000000000000000000111100000000000000000000000000000000010000100111011111111101000000000000001111111101100000000011011110000001010111101111111000101111010000000000000000000101111000000000000000000000000000000010111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                 
    249: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011001001111000001111000111111000000000000010001100001111111111100000000000000000010000000000000111111111110110111101111111101000000000000000000111110000000000000000000001000000000000110110111111111010000000000000000001111111110100000001011111111000000111110110111101000111111100000000000000000000011110000000000000000000001001000000011111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    250: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000000000000000000000000000000000000000000111000001111000001101000111111000000000001001000100000111111110110000000000000000000000000000011011110111111110110111111111110010000000000000000111010000000000000000000000000000000101011111111111010010000000000000000001111111110110000000011101111100001111111111111110101111111000001000000000000000011110000000000000000000000000101010001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    251: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001111000001000000000000000000000000000000000000000101100011101000001110000111010000000000000110000100000111111111101000000000000000000000000001101111011111111000011110010111111100000100000000000111100000000010000000000000010101111111111111111100100000000000000000000011111111101000000000111111111010000111111111111111001111110000100000000000000000111110000000000000000000000001101010101111111100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    252: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000011110000000000000000000000000000000000000000000000111100000111100000111000011111100000000000010001110000011110111111110000000000000000000000110111111111110011101111101001111111010000000010000010111110000000000010000000010101011111111111111010010000000000000000000000001110111110101000000011111111110000011111111111111111111111000000000000000000000001110000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                 
    253: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000111110001111000000111100011111100000000000001000111000011011111111111101000000000000000010111111111111001100101100100101111111111000000000000000111111000000000000001101011111101111110111010000000000000000000000000000011111101110100000000001111011111001011111111111111101111100000000000000000000001111011000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    254: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100000000000000111101000000000000000000000000000000000000000000000111100100111100000110100011111100000000000011000001001001000111111110110100010000010101111111111111101010111110100000111011111111100000000000000111110100000000011101111111111111110111000000000000000000000000000000000011111111100110000000111101111101000101111111011111111101100000000000000010000000111100000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    255: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001011100000000000000000000000000000000000000000000000011100001111000000011000001111110000000000000100110000001001011111111111111000101010111111111111111100011111111000011101111111111011010001000000111111001011111111111111110111110101000000000000000000000000000000000100101111111110101000001011100011110000011111001111011110111000000000000000000000000111100000000000000000000000011111100111101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    256: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000111110000111100000011110001111101000000000010100001000000100110010111111111111111111111101111111110001111110110000101010101010111111111111010001011111111111111111111111111111100000000000000000000000000000000000000000111111111100010000000011000111111000111111111111111111111100000000000000000000000101110000000000000000000000111110110010111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    257: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000111101000111100000011000000111110100000000000110001100000110011011111111111111111111111110110111100001111110010001110011100001111111111101111111111011111111111101111111111110100000000000000000000000000000000000000000111111101110110000000011000011111100011101000111111111110000000001000000000000000111100000000000000000000000011111100000010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    258: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000111110001111010000011110001011111000000000000001000100000001010010110101111111111111101010111111100111101110010110001110000011111111111111111111111111111011111111011111111111110000000000000000000000100000000000000011011111110110110000000111100011111100011111000011111111111100000000000000000000011111010000000000000000000001111111000000000101111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    259: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000000000000000000000000000000001000000000000001111110000101100000001010000111111110000000000000001100000000110001011011010110001010000001111100001010111000000100101100010110110111111111010011111111111111111111111101111011110000000000000000010010000000000000000101111101100100101000000110000111111101011111100000111111111111000000000000000000000111100000000000000000000000111110100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    260: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101000000100010000000000000000001000100000000000000111101010111100000000000000111111010000000000000000110100000010011011000101010100000000111111010001111010100001010111001001111001001010100001001110110111011011111111111111111111100001000000000000000000000000100000111111111010100110000010011000011111110001111100000010111111111111110100000000000001111000000000000000000000001111111000000000000110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    261: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000001101001000000000111110000111100000000000000011111110100000000000000010000000010001011011001110000000011111111000111110110001011000110001110100000111100000000011110011011001110111111111111111111111000010000000000000000010000000010111110001101100110000000111000001111111011111100000011111011111111010000000000000001111100000000000000000000001011111000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    262: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000111100000000000000000000000000000000000100000000000001111111000111100000001000000011111111000000000000000011000000000010011001000000000010111011100011111011010000101011010010110000111000000000000001110011011000111111111111111111111111101000000000000000000000000000011111110100001100110000000011000110111111111111100000001111101010111010000000000000010110000000000000000000000001111110000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    263: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100100000000000000000000000000000000000000000000001111110001111100010000000000011111110100000000000000010100000000011010101000100000101101110101011110011000001100010001111000011010000000000000011100001001100101011111011111011011111111010100000000000000000000011111111010011001100110000000110000011111111101111100000111110000001001000001000000001011111000000000000000000000001110111000000000100010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    264: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110101111000000000000000000000000000000010000000000100111111100011110000011101000000111111100000000000000001010000000000010000000000011111000011000101111101000001000101010100000101101000000000000001110001010010011111101110101111101011111111101000000000000000000010111111000111000101010000000111000001111111111101111000010101000000000000000000100000101111000100000000000000000001111110100000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    265: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111110111000000000000000000000000000000000000000000001111111001111100000001110000001111111110000000000000000110000000001000000000001011100111001011110110110000101011100110100000110000000000000000001110001010111001011111011101011101011111111111100000000000000101011111111100010010100111000000011000011011111111111100000011100000000000000000000000000011111000000000000000000000011111110000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    266: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110011111100000000000010000000000000000000000000000001111111000111100000001111100001111111100000000000000000011000000000000000000101010100011001111011011010000101010101110000010100000000000000000001100000010001001111111011110001110001011111111110100000000100111111011100001100011000000000001011000011111111111111110001111110000000000000000000000000111101000000000000000000000001111111000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    267: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000010001000000100000000100000000000000011111111100011110000001111100000111101110100000000000000100000010000000000000001000011100010100011101000000010111010100000101010000000000000000101110000100010100110111000111100111001111111011111010010110111111111111100000010001100100101000110000011111101111111111000111000000000000000000000000000111110000000000000000000000011111100000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    268: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110001111110000000000000000001000000000000100000000000110111100101111000000111111000111111110000000000000000011100000000000000000000100101010111010101111000001010100011000100011000000000000000000010110000000000110011101100010100001100001011111111111111111111111111110110000000010000010000000011000001111111111011011000111100000000000000000000000000101111000000000000000000000011111111000000000000101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    269: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110010111100000000000000000000110000000000100000000011111111100000111100100111101000011111111000000000000000001010000000000000000000000100011011000111110000001011100110000001100000000000000000000001010000000000000000111110000111001111001011111111111111111111111101111001000000001000000010000111000011011111111111111101110000000000000000000000000000111110000000000000000000000011111110000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    270: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111000001110010000000000000000100010000101000010000000011111111100000111110000111100001111111111001000000100000000100000000000000000000011000011000011111100000000000010010000001110000000001000000000011110000000000000000110101000101000001000001011101111101111111011100110000000000000000000010000011000011111110111111111110111000000000000000000000000001111010000000000000000000000001111110000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    271: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000111110000011000000000000000000001010000000000000000000011110110100001011110100111110000011111111100000000000000000010000001000000000000000101110000001110100000000100011000000010000000000000000000000001010000000000000000110111010011100001110000001111111111111110101101010000000000000000000101000111000011111011111111111011110000000000000000000000000001101110001000000000000000000011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    272: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000100000001100001000101000000001111111110000001111010011100000111011111000000000000000000000000000000000000000000011000000111111000000000000101000000011000000000000000000000001110000000010000000011001100000010000011100000001101111111011001011100000000000000000000010000101000001111111111111111111110000000000000000000000000101111110000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    273: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000001010000100100100010011111111110000001111101011010000011111111100000000000000000000000000000000000000010111000000111110000000000000100000000011000000000000000000000000010000000000000000011100110000011000001110000000111110101100011101000000000000000000001010000011000101111111111110111111010000000000000000000000000011111110000000000000000000000001111111000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    274: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000010000000110010100000000001011111111110000000111110111000000111101111110000000000000000100000000000000000000010000000010101010000000000000100010001100000100000000000000000000000000000000000000001010011010001100000111000000001011000110011110000000000000000000000110001101000111111011011111111111100000000000000000000000000011111110000000000000000000000011011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    275: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010000000000000000000000000100001011000010010100000101111111100000001111100011000000011111111101000000000000000000000000000010000010101000000011010100000000000010100000000100000000000000000000000000000000000000000000001100000000000111000001110000000000101100011100000000000000000000001100000110000011111001111111101111111100000000000000000000000011111110000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    276: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000001000001000000001000000111111111111000000111110110100000011111111110000000000000000000000000000000001000100000000101101000000000000001000000000110000000000000000000000000000000000000000000000111000000100010100000101000000101100100111000000000000000000000000111011110000011111000111111011111110111100100000000000000000011111101000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    277: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000010000001010011000100000011110111111000000011110010100000011111111110100000000000000000000000000000000010000000000010010000000000000010000000001000000000000000000000000000000000000000000000000010100000000010110000000000000000000000001000000000000000000000010100001110001011111001011111001111111111110100000000000000001011111110000000000000000000000001110111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    278: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000001000001010000100100000111111011101000000111111111000000011111111111000000000000000000000000000000000000000000001010100100000000000101000000011000000000000000000000000000000100000000000000000011000000000000110000010000000000000100000000000100000010000000011100010100001111111001111111001111111111111100000000000000001111111111000100000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    279: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000110000101001000000001110111111110100000011110010000000101110111110100000000000000000000000000000000000000000000001010000000000000100000000000010000000000000000000000000000000000000000000000001110000000000011100000000000000000000000010000000000000000000001100001000000111111000111111001010010111111010000000000000001011011110000000000000000000000001111111000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    280: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000010100010000010011000111110111111000000001111011100000011111001111100000000000000000000000000000000000000000000000000000001000001010000001001000000000000000000000000000000000000000000000000000101000000000001010000000000000000000000000000000000000000000111001000000001110111001101111001111001010010000000000000000001111110111100000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    281: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000010001101001000000111110011111100000011111011010000011111011111110000000000000000000000000000000000000000000000000000000000000100000000100000000010000000000000000000000000100000000000000000110100000000000111000000000000000000000000000000000000000000111100000000001111101001111011001100000001000000000000000000001111110011100000000000000000000001111111100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    282: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000010100010100100101001111110111110010000001111101000000011111011111100000000000000000000000000000001000000100000000000010000000010000000000010000000000000000000000000100000000000000000000001000011000100000000001100000000100000000000000000000000000000000110000000000011111100001111110011100000000000000000000000000111111000010101000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    283: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010000000000000000000000000001000000010000100110010001111100011111000000011111101000001111111101110111000000000000000000000000000000000010000001000000001100000001100000000000000000000000001000000000000100000000000000000000000001110000000000000110000000000000000000000000000000000000011111000000000011100010010111111011010000000000000000000000000011111100011110000000000000000000001110111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                  
    284: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000101000010000010010111110101111100000001111110000000011111010111110100000000000000000000000000000000000000000000000010010000010000000000000000000000000000000000010011010100000000010000000000000110000000000000001000000000000000000000000000000000000001110100110000011110000001111110111000000000000000000100000000111111101001111000000000000000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                   
    285: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001100011011011001111110010110100000000111011000000111111001111110100000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000011111111110101000001000000000000011100000000000001000000000000000000000000000000010000011110000100100011110000011111111111000000000000000000000000000010110000111111110001000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                   
    286: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111000000000000000000000000000000000000000110001001001011111010011111100000001111100000000111111101111111010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001011111111111000000000000000000000001110000000000000000000000000000000000000000000000001011110000110000011110000001111111100000000000000000000000000101111111001111011101000000000000000000011101111000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                   
    287: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000001000000000000000000000000000000001010010100101001101100011111010000001111110010001111111010111111100010000100000000000000000000000000100000000000000000000000000000000000000000000000000001010111111110111110000000000000000000000111000000000000000000000000000000000000000000000010111110111110000111110000111101111110000000000000000000000010011111110001101100111000001000000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                   
    288: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111010000000000000000000000000000000000000001001010101111111110011111100000000111111000011101111101111111110000000000000000000000000000000000011000000000000000000000000000000000000000000000000000011111110111111111110000000000000000010001110001000000000000000000000000000000000000000001111110001111100011110000011111111100000000000000000000000000001111111110110001111110100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                   
    289: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000111101000000000000000000000000000000000000000101001110110011111100011111110001000111101000011111111100111111111000000000000000000000000000000001010000000000000000000000000000000000000000000000000001111111111111111111010000000000000000000001011000000000000000000000000000000000000000000111111110111111000001010000011110111001000000000100000000000000111110111111110000111111010000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                                   
    290: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000001100101111101111100001111000000010111110001101111111111111111111100000000000000000000000000000000000100000000000000000000000000000000000000000000100011111111111111111111111000000000000000000000111100100010000000000000000000000000000000000111110100110111100011100001011111111000000000000000000000000000111110011111000011111011111010001000000010111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    291: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001111110000000000000000000000000000000000000000000000110111111111000011111110000000111111000111011101001111111111010000001000000000000000000000000010000000000000000000000000000000000000000000000001110111011111111111111111110000000000000000000001010000000000000000000000000000000000000011111011100111111000011110100111111100000000000000000000000000011111101011111110011100001111100000000000000111111110000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    292: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000100000000110011011111111100001111100000000011111011010101111110110111111110000000000000000000000000000000000000000000000000000001000000000000000001000000001011111111111111111111111111100000000000000000000011101000000000000000000000000000000000001111111010011111100001100001111111110000000000000000000000000000111100000111100111110001111111000000000000010111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    293: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000011011101110111100001011110000000111111001100111111101111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111010110111111110110000000000000000000000101010000000000000000000000000000000011111101100111111100001110001111111100000000000000000000000000011111100100011010011000000111111000000000000011011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    294: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000001101111111111000001111010000100011111000100111111101110101011111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111101111111111101111111111000000000000000000000000001000000000000000000000000000001101101101100111110100101110010111111100000000000000000000010001011111000000111111111100011111111000000000000001111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    295: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000001011111111111100011111100000000111111000000011111100111110111111110000000010000000000000000000000000000000000000000000000000000000000000001010111111110111111111111111110111111110000000000000000000000000000000000000000000000001000000111110111100111111000001100011111110000000000000000000010000000111110000000001111111000111111011000000000000000101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    296: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101000000000000000000000000000000000000000000000111111111111000000111111000000011101100100011111110101001011011111100100000000000000000000000000000000000000000000000000000100000000000000111111111111111111111111111111111111111010000000000000000100000000000000000000000000000000011010100001010010111100001111111110111000000000000000000000000011111111000000000011111110101101111100000000000000011111111000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    297: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011110100000000000000000000000000000000000000000000011111101111000010111100000000011110100000001111110111110011111111100000000000000000000000000000000000001000000000000000000000000000000000011011101111110111111111111111111111111101000000001000000000000000000000000000000000000000011100110001101111111100001110011111111000000000000000000000000001110110000000001000111111111010111100001000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    298: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000010101111111011000001111110000000011111100000111101100101010011111111110000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111111111111011111111100000000000000000000000000000000001000000000000010100000101100111111000001111111111101000000000000000000000000111111110000000000010011111111111110000000000000000010011011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    299: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001000000000000000000000000000000000000010000011111111111000001111110100000011111000000001111110010110011011101111000010000000000000000000000000000000000000000000000000000010000100011111111111111111111111011111111111111111111010100000000000000000000000000000000000000000000101000000010101111111100000111111111100000000000000000000000000011111000000000000000101011111101111010000000000000000101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    300: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111000000000000000000000000000000000000000000000001111111111000000111111000000001111110000001111100101101001101111111100000000000000000000000000000000000000000000000000000000000000011111111111110101111111111111010110101101101101111000000000000000010000000000000000000000000001010000000001000011101100001011111111110000100000000000000000000111111100000000000000000001011111100000000000000000000010111111110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    301: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000001011111111000001011101000000001111011000001111110000101000001110111110000000000000000000000000000000000000000000000000000000000000001111111010000000001111111001111011010101010111111110000000000000000000100000000000000000000000110000000000001111111000000101111011100000000000000000000000010111111100100000000000001000001010000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    302: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110111000000000000000000000000000000000000000000000001111111110000001111111000000001111100010001111100011101011001111101110000010000000000000000000000000000000000000000000000000000000111111111010000000000110101000000000000000000000111111100000000000000000000000000000000000000000100000000000000111111100000010111111100000000000000000000000010111110000000000000000000000000000000000000000000000000000001111111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    303: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000000000000000000000000000000000000000000001111111010000000111111000000000111111000001111110001010001001111111111000000000000000000000000000000000000000000000000000000000011111111100000010000000001000000000000000000000000001111111000000000000000000000000000000000000001000000000000001111111000000001111111110000000000000000000000011101111000000000000000000000000000000000000000100000000000001011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    304: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000011111110000001111111110000000111111000000111110101101001100111111110110000000000000000000000000000000000000000000000000000000011111101010000000000100000000000000000000000000000000111110110010000000000000000000000000000000000100000000000000111111100000000111111100000000000000000000000011111100000000000000000000000000000000000000000000000000000000001111111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    305: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101000000000000000000000000000000000000000000000101111101000000111111100000000011111110001111110000110100001111111111010000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000001000001111111000000000000000000000000000000000010001000000000000101111100000000111111110000000000000000010000001111110000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    306: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000111111100000000111111110000000011111111101011110000010011001111011111110000000000000000000000000000000000000000000000000100010111111100000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000011111111100000000111011100000000000000000000000111111000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    307: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011111000000000000000000000000000000000000000000000000010111100000001011111100000000001101111111111111100011001000111001111111000000000000000000000000000000000000000000000000000111111010000000000000000000000000000000000000000000000000000001111101100000000000000000000000000000000000000000000000111111000000000101111101000001000000000000000111111100000000000000000000000000000000000000000000000100000000000001111111101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    308: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000011111100000000111101111000000000111111111111111110010001001011001111111100000000000000000000000000000000000000000000000001111111110000000000000000001000000000000000000000000000000000000011111010100000000100000000000000000000000000010000000110111110000000111111110000000000010000000000111110000000000000000000000000000000000000000000010110101100100000000101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    309: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111000000000000000000000000000000000000000000000000001101110000000111111111000000000011111111110111000010101001111001101111101000000000000000000000000000000000000000000000010111111010000000000000000000000000000000000000000000000000000000011111110000000000000000010000000000000000000000000000111111100000000111111101000000000000000000000101111000000000000000000000000000000000000000000011111110111011001000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    310: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001111111101101000000000000000000000000000000000000000000000101111100000001011111111000100000001011111111111100010011001111001111111110010000000000000000000000010000000000010000001111111110000000000000000000000000000000000000000000000000000000000001111111100000000000000000000010000000000000000100000011110110000010111111110000000000000000000001111100000001000000000000000000000000000000000000111111111111101101111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    311: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111011011100000000000000000000000000000000000000000000000011111110000000111111101100000000010100101111110000001001100111000110111111100000000000000000000010100000000000000000000111111101001001000000000000000000000000000000000000000000000000000001111111000000000000010000010000000000000000000110000011111100000001111111100000000000000000010011111100100000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    312: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111100110000000000000000000000000000000000000000010000001111100000001111111111100000000000010001111111100000011000101101111111111000000000000000001000001010000001000000000000111110100000000000000000000000000000000000000000000000000000000000000111111111010000000000000000000000000000000000110000101111100000011110111100000000000000000000001111110000000000000000000000000000000000000000000000111111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    313: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000110000000000000000000000000000000000000000000000000111101000000111011111110000000000000000111111100000001100011000010111111110100000000000000000101100000000000000000001111111000000000000000000000000000000000000000000000000000000000000000011111110000000000011100000000000000000000000110000101111110001011111011110000000000000000000011111111000000000000000000000000000000000000000000000011110111111110111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    314: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000111000000000000000000000000000000000000000001000011011110000001111111111111000000000000000011111110000010010001011010111111110000100000000000000110100000000000000000101111101000000000000000000000000000000000000000000000000000000000000001100110111000000010001100000000000000000000101110000101111100000011111110000000000000000000001011011110100000000000000000000000000000000000000000000001111110100111011011111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    315: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000110000001000000000000000000000000000010000110000001111100000000111111111110000000000000000101111110000001000011001101111111110000000000000000000111000000000000000100011111100000000000000000000000000000000000000000000000000000000010000000111011011010010000001110000000100000100000011100000011111100000111111110000000000000000000001111111111010000000000000000000000000000000000000000000000111111110000101100101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    316: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011101001011000000000000000000000000000000000000001111110000111111000001111111111111100000000000000001111111000011100011000010111111111000000000000000001110000000000000000000101111000000000000000000000000000000000000000000000000000000000000000000100111001100000000000011000000000000000000101111000011111110000111111101000000000000000000000111111111101000000000000000000000000000000000000000100000011111111000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    317: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000011100000000000000000000000000000000000001010111000111111000000110111111111110000000000000001011111100001000011010101010111111000000000000000010110001000000000000000110111000000000000000000000000000000000000000000000000000000000000000000100001000110000000000011000000000000000000001100000011111100101111111100000000000000000000011111111111110100000000000000000000000000000000000000000000000011111110000000000011111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    318: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000101000000000000000000000000000000000000001110101000111111000010111101111111110000000010000000111111000001000001001001111111111000000000000000111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000110100100000000000001100000000000000000011110000011101110011111111000000000000100000001011111011111111100100000000000000000000000000000000000000000001011111110000000000011111111100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    319: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000011100000000000000000000000000000000000000100011101011110001001111111110111110100000000000000011101110001000011000100101011111100000000000100111100000000000000000010111110000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001010000000000010000101110001011111100101111100100000000000000000001111111101111111110000000000000000000000000000000000000000000000011111111100000001000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    320: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110110000001010000000100000000000000000000000000001110011100111111000000111111111111111000010000000000001111110000000001100101010111110100000000000001011000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001010000001011111000101111111111111110000000010000000000010110111001111111101000000100000000000000000000000000000000000000000111111101000000000011110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    321: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000001110000000000000000000000000000000000000111101110011111000000011101111111111100000000000000001111111000000010100000110111111110001000000001110000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001010000001110111000111111111111111110000000000000000000011111101000011111111100000000000000000000000000000000000000000000000011111110100000000000111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    322: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000110100000000000000000000000000000000000001110001111111100000001111111101111110000000000010001111101000000001011100010101110100000000000001110000000000000000000001110000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001110000001111011000011111111101111101001000000000001000011111100001111111111000000000000000000000000000000000000000000000000001111111000000000001011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    323: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111000000000110000000000000000000000100000000000000000001010111111000000011111110111111111000000000000000111111100000001000001101110111110000000000011100000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100010100000010111111000111111011111101100000000000000000000111111100000011111111110000000000000000000000000000000000000000000000000111111100000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    324: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000010000001000000000000000000000000000000011000000000011111110000000000111111111111101100000000000000011111100000001001100100010111110000000000011100000000000000000000001100000000000000000000000000000000000000000000000000000100000000000000000000010000000000000000000001010001111000011111111000011111111110111110000000000000000001111110100000011011101110000000000000000000000000000000000000000000000000011111110000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    325: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000010100000000000000000000000000100000100000000011111111000000000011111111111111110000000000000101110110000001000100010100111110000000000010100000000000000000001001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001110000011111111100111011111111101110000000000000000001111111000000011111111101000000100000000000000000000000000000000000000000001111111000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    326: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000000000000000000000000000000000000000100000100001111111100000000000011111111111111111000000000000111111110000001001101100100111111000000001010000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011001110000101111110000111111101100101110000000000000000111111111000000011111111110010000000000000000000000000000000000000000000000000111111100000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    327: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101110000000000000000000000000000000000000100000001000000011111101101000000000001111111011111110100000000000001111100000001100100110100111110000000000110000000000000000000000010100000000000000000000000000010000000001000000001000000000000000000000000000000000010000000000000000101000101000111111011001011110111011101100000000000000000101110110000000001111111111000000000000000000000000000000000100000000000000010111111100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    328: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000100000000000000000000000000000000000000010111111000000000000100110111111101111001000000000001111111000000000100010110011111101000001110000100000000000000000011000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001100000000111111111000111111110110101110000000000000010111111111000000011111111111100000000000000000000000000000000000000000000000000001111111000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    329: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000001111011111000000000000000111111111111111100100000000100111110100000100110101010111111000000000101000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000110000001011111110000111111111000101010000000000000011111111111000000001101111111100000000000000000000000000000000000000000000000000101111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    330: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010000000000000000000000000000000000000000000000000001111111000000001000000000011111111110111100010000000001111111000000001001010100111111000000001100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100110000001001111110000111111111010011100000000000000011111111100000000001111011101100000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    331: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000111111101000000000000000000101111111111110110000000000001011111000000000100101010111011100000011100000000000000000000000010000000000000000000000000000000000000000001010001010000000000000000000000000000000000000000000000100001010000101101111110000111111111001011110000010000000101111111111000000001111111111110000000000000000000000000000000000000000000000000010111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    332: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011111110100000000000000000000000000000000000000000000010101111110000000000000000000001101111111111101000000000000111111110000000100010100111111110100001100000000000000000000000000000000000000000000000000000000000000000000100000000000010010000000000000000000000000000000000000010000111100000010111010000011111111010000100000000000010111111111110000000011111111111111000000010000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    333: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001011100000000000000001000000000000000000000000000001011111111000000000000000000000000111011111110110000000000000111111000000000101010110011111100000011100000010000000000000000000000000000000000000000000000000000000100000010000100000000000000000000000000000000000000000000000010000001000000001111111001011011111001001110000001000011110110111110000000001111111111101000000001000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    334: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000001111110111000100000000000000000001011110111111111100000000000111111110000010000110101111101100000011000000000000000000000000000000000000000000000000000000000000000100001001000100000000000000000000000000000000000000000000000011000011100000011111000000111111011101011000000000000011111111111111000000001111111111111000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    335: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000111111111110100000000000000000000000011111111111111010000100000011111100000000100101010011111110000011000000000000000000000000000000000000000000000000000000000000000100000100001010000110000100000000000000000000000000100000000001000001010000010111000000011111111001001110000000000111111111111110000000010111101111110100000000000000100000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    336: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000001000001111111111000000100000000000000000011111111111111101000000001011111110000000001010100101111111000011100000000000000000000000000000000000000000000000000000000010010010000100000110000011100000010000000000000000000000000000000010100001100000011111000000111111110110001000000000001011111111101111000000001110111011111100000000000000000000000000000000000000000000000000001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    337: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000010111011111111000000000000000000000000000111111011111111100000000001111010000000000011010010110110000011000000000000000000000000000001000000000000000100000000000000000100000010001010001011010100000010000000000000000000001000000001100000101000010111000000011111111001100100000000011111111001111111000000001111001111111100000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    338: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101110000000000000000000000000000000000000000000011111111110111000000000000000000000000001101111111111111111000000011111110000000001001010010111111001011000000000000000000000000000000000000000000000000000000000001000100000101101111001111001100000000000000000000000000000000000000110000110001011000000000110111101100011000000000011110101011111011000000101110000011111110000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    339: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000001101111110111111000000000000000000000000000011111111111111111100000011111110000000000110100001111110000110000000000000000000000000000000000000000000000000000100000001000110001111111111111111110110000000000000000000100000000010000000101000111000101001000000011111110111010000000001111011100011101110000000011110000111111100000000000000000000000000000000000000000000000000000001111110000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    340: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110001000000000000000000000000000000010000011111111111011110100000000000000000000000000011111111110111111010000001111110000001000010010100111111000111000000000000000000000000000000000000000000000000000000000010101000011110111111111011111010100000000000000000000000001000000000010000001000000000000000111111101000011010000000111111110001111111000000101110000001111111100000000000000000000000000000000000000000000000000010111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    341: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000101111111111111101111100000000010000000000000000001111011111011111101000001111111000000000011000000111111100010000000000000000000000000000000000000000000000000000000100001000110101111110111111111111110100001000000000000000000000100000000011000011100000000000000011011101111011000000011111111100001111111100000011000000001111110100000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    342: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111110000000000000000000000000000000000000111111111011100001111000000000000000000000000000000111111111111111101000001111110000000000010100000110110101101000000000000000000000000000000000010000000000000000000010001001111111111111000111011111111110000010000010000001010000100000000001000001000000000000001111111100100001001001111111111010011111111000000101010000000111111101000000000000000000000000000000000000000000000000010111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    343: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000001000000000000000001011011111111010001111100100000000000000000000000011111111111110111111110001101110000000000001000000011111000110000000000000000000000000000000000000000000000000000011011001000111111111000010000001111111111000000000000011100000010100000000011000011000000000000000111110001011000000000101111011000000111111000000001000000001111111110000000000000000000000000000000000000000000000000000101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    344: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110000000000000000000000000000000100111111110111111000000011010000000000000000000000100011101111111111101111111000111111100000000100000000111111101100000000000000000000000000000000000000000000000000000001010010111111111100100000000100010111111100000001001101110110001010000000001100001110000000000000011111100001000000011111101111000001111111100000000000000000111111101000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    345: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000010010000011111111111111111000000111100000000000000001000000001011010111110110000110111101111110000000000000000000011110101100000000000000000000000000000000000000000000001000000001001001111111110100000000000000010101111111000001111111111111000011000000001100000100000000100001111110001001000000011111110111000000110111100000000000000000101111111010000000000000000000000000000000000000000000000000011111010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    346: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111010000000000000000000000000000001011111111111011100000010011100000000000010000000000001110001011111111000111010000111111000000000010000000011111001100000000000000000000000000000000000000000000000000000011001111111111010000000000000000000011011111110101111111110110000001000000000100011110000000000001111110000001000000011110101110000000111111100000000000000000111111111100100000000000000000000000000000000000000000000000010111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    347: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110100000000000000000000000000000101111010111111111110010000011110000000000000000000000111110000111111111000000101001111111000000000000000000101111101100000000000000000000000000000000000000000000000000000010111110111101100000000000000000000000111111111111111111011111100110000000000100000100000000000001111010000000000000110101001110000001111111010000001000100000011111111110000001000000000000000100000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    348: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000001111111100011111111000000000001010000000000000000000010011111100111111111100010000000011111000000000000000000011110101000000000000000000100000000000000000000001000000000000011101111111110000000000000000000000000001011011111111010111111100000100000000110001010000000000001111100000010000101101010101011000000011111100000010010000000001111111111100000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    349: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110001000000001000000000000000111111000001011111111100000000000101000000000000000000001111111110111101111110000000000101111100000000000000000001111101100000000000000000000001000000000000000000000000000000010111111101110000000000000000000000000001011111111101000001111110010000000000010000101000000000110111110000000100000110100010110000000101111110000011011000000010111111111110000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
    350: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101110000000000000000000000000111101101000101111111110000000000000100000000000000000000001010111111011111111100000000100111111010000000000010000001111111000000000000000000000000010000100000000000000000100000011111111110000000000000000000010100000000000110100100000000111100001100000000100000100000000000011111000000000101000000011000010000000111111100000011111100000001110111111111000000000000000000000000000000000000000000000010111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                      
    351: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000000000000000000101011110000000011110111010000000000000000000000000000000000011110000111111111111110000010000111111100000000000000000001111110100000000000000000000000001000000000000000000000001011111111111101000000000000000001001100000000010000010000000000111110000010000000110001110000000000111111000000001000000000100011100000000011110100000111011100000011111101111111110010000000000000000000000000000000000000000001111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                      
    352: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011000001000000000000100011111010000000111111111110000000000000000100000000000000000101110000011111111111111000000000101111000000000000000000001111111000000000000000000000000100100000000000000000010100101111111110100000001000000000000011101000001000100000101000000001111010100000000010000010000010001111111000000010100000000000000100000000001111110000001110110000000111001011111111000000010000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                      
    353: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110100000000000000000011111100000000010111011111110000000000000000000000000000000000111111010001111110111111100000000111111100000010000000000000110110001000000000000000000000010010000000000001111111111111110110100000000000100000000001001100100001111111000100000000001111000100000000011000101000000001111101000000100000000000000000100000001011111110000000111110000001111101111110111110000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                      
    354: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000001111000000000000011111011111000000000000000000000000000000000000111011110001110111111110000000000011111100000000000000000001111110000000000000000000000001001000000000101110111011111111111010000000000000001000000101101111001111111111100111000000000111000110000000010000110000000010111101000010100000000000000000000000000010111110000000010000000000111000011111111111000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                      
    355: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000100000000000111110101111100000000000011100000000000000000001011111111110111111101111100000000011101101000000100000000000111110000000010000000000000000100010000010011111111111111110101000000000000100100000010000111110001110100011110001100100000111100010000000011001010000000011111100000010000000000000000000000000000011111100000001001000000001111000011111110111110001000000000100000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                      
    356: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000001111110011110000000000000010111001000000000000001110101111111111111111111110000000001111100000000100000000001011110000000000000000000000011001000100001111111111111110100000000000000000011010100000000101111011110000001110011110010100001110101000000010000100000000111111100000100000000000000000000000000000011111111000000000000000000101100001111111011011000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                      
    357: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000100000010111100011111000000000000011111000000000000000001110000001111111111111111110000000101111110000000010000000000011110000000000000000000000001001000010111111111111100000000000000100000000101010000000000101111101110000000111001100111100011110111000000011000110000010111110100100000000000000000000000000000000011111110000000000000000000111100001111111101111110001000000000000000000000000000000000011101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                      
    358: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011011100000000000000000000000000100011011100011111000000000000001111000000000000000001111000101111111111111111110100000011111100000001000000000001011110000000000000000000000100100000001111111110000000000100000000111000000011011100011101111010111000000000111110100110100001110101000000011000100000011111110000000100000000000000000000010000000011111010000000000000000000110100001011111100111011000000000000000000000000000000000100011111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;                      
    359: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000001111010100111110000000000000010111000000000000000101111111111011111011111110111000000001111110000001101000000000111100000000000000000001000100010000011111111110100000100000000011111111000001100000001111111111111000000000111011101111110010111111000000011001110000011110110000000000000010000000000000000000000011111100100000000001000001011000000111111110001111100000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;                     
    360: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000100111000011010010000000000000111010000000000000011111111011111101111111011111000000001111111000000100000000000011011000000000000000000001101100001111101111000000000000000000010111111000011110100111111111111011100000000011111110111111101111111100000011000000000101111010000000000000000000000000000000000001011111110000000000000000000111100000111111111001110111100000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;                     
    361: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111101000000000000000000000000011101111000111110000000000000000001000000000000000011010111111111000110111101111100000000111110100000100000000000111100000000000000000000000100010000111110111000000000000000000011101011110001111000011010111111110100000000001111111110111111101010100000011101110001111111100000000000000000000000000000000000000001011100000000000000000000011010000011111111100011101010000010000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;                     
    362: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110100000000000000000000000100101100000111100000000000000000000000000000000000111000011011111000111111000111110000010111110000001110000000000011100000000000000000000010011000011111111101000000000100000000011100011100010110010111010111111110100010000011111111100011011111111000000110101000001111111000000000000000000000000000000000000000111111110000000000000000001111000000110111111101000101011000000000000000000000000000000011101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    363: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001111111000010000010000000000001100011110000111010000000000000000000000000000000010111000000111110100111110100011110000000111111000000100000000000111110000000000000000000111000001111111111000000000111011000000011000101111001111001110000011111110000000000001011111010011111001111100000011001110111111110100000000000000000000000000000000000000111111100000000000000000000010000000011111111110010100101010000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    364: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011110000000000000000000000001010111110001111100000000000000000000000000000000000101000000011110000011111000001111010001011011000001010000000000111100000000000100000000000011000101111111000000001011111101000111100000110011111000111000011111111000000000001111110000001111000111100000111111000001111110000000000000000000000000000000000000000111111100000000000000000000101000000011111011101000110010101000000000000000000000000000101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    365: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000001000110100000111100000000000000000000001000000000001110100100001110000011111100000011000000111111100001010000000000011110000000000000100000111000011110111100000000001111111101000011000000111001110011100000000111101000000000001111110000001111010111100000011011101111111100000000000000000000000000000000000000001011111100000000000000000000100000100011111101101100011000000100100000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    366: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111000000000000010000000101001111100001111010000000000000000000000000000000000110110111111110000001111100000001100000111110100001010000000000111000000000000000000101000100011111110100000000011111111111001111000000011111110101100000011111110000000000000111000000001111001111100000111110011101011100000000000000000000000000000000000000001111111100000000000000000000000000000011111111100100001100100100000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    367: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000001000110011101000000111100000000000000000000000000000000001111111111111110000011111110000000110000011111000000100000000000011110000000000000000000101001111111110000100101110110101111000111000000011101111011100010001111110000000000001111100000001111000111010000111111101111110000000001000000000000000000000000000000000111111000000000000000010000000000000001111101100110000110000010000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    368: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111000000000000000000010100010001000001111000000000000000000000000000000000000111111110110110100000111111000000001100010111100001110000000000111100000000000000000011110100111111101000001010111110010111101101010000001111111111000000010111111000000000001101000000010111101111100000011111011111111000000000000000000000000000000000000000011111111100000000000000000000000000000011111100110001000001000000000000010000000000000000010111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    369: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000001100011000100001111100000000000000000000000000000000000111000000111110000001011111110000010100011111100000110000000000011110000000000000000001010011111111100000011111111010000011111110000000001111111111100000001011100000000000001111000000001111100111100010111101111111110010000000000000000000000000000000000000001110111000001000000000000000000000000001111100111011100001100000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    370: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000010000101010000001110100000000000000000000000000000000010110100000011100000000111111010000001010001111100000110010000001101100000000000000000101110011111111000011111111100000000101111110000000000111111110000000001111110000000000011101000000011110100111100000111110111111000000000000000000000000000000000000000000011111101000000000000000000000000000000011111100010000110000110000000000000000000000000000001011110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    371: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011011100000000000000000101000100101000101111000000000000000000000000000000000001111000000001110000000011101110000000100011111110001100100000000111010000000000000000011011111111100001111110010110000000111111100000000000111111111000000000111010000010000011110000000011111001111000001111111111111000000000000000000000000000000000000000000011111110000000000000000000000000000000011101100110001010000101000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    372: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000110000000110000011111100000000000000000000000000000000000011101000011100000000001111111100000000000111110000110010000000111100000000000101000111100111111101000111010001110000000011111110000000000011111100000000000111100000000000101100000000010111110111100001111111111110000000000000000000000000000000000000000000101111110000000000000000000000000000000001111100001000011000001000100000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    373: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000001000000100010000001110100010000000000000000000000000000000011110111111100000000001111111010000000001111111000111010000001000000010000010100000111111101101100111111000001111000000011011000000000000101111110000000000111100000000000111110010001111111010111100000111111101110000000000000000000000000000000000000000000111111101000000000000000000000000000000101111010101000001000001100000000000000000000000000001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    374: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110100000000000000011100000001100000011111010000000000000000000000000000000000011111011110000000000000111111100000000000110111000100010010001100000000000001000001111111111110000011110000000111000000011111100000000000110111100000000000111100000000001011001011101111110001011100111110111111100000000000000000000000000000000000000000011110111000000000000000000000000000000000011111100010100011100000100000000000000000000000000001111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    375: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000101000000010010000011111000000000000000000000000000000000000000111111010100000000000010111111000100000111110001111110000000100000000100011100000111111111111001111000000000111100000111110000000000000011111100000000010111010000000011111111101111111111101111000001111111110000000000000000000000000000000000000000000001011111100000000000000000000000000000000011111000001000001100000011000000000000000000000000010111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    376: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000010000000001100000001111100000000000000000000000000000000000000010101000000000000000001111111000000000011111100110011000001110000000000110000101111111111100011101100000001011010000011111100000000000011111010000000000111111010000111111111111111101111000101000011111111111100100000000000000000000000000000000000010011111110000000000000000000000000000000000010111100000100000101000000000000000100000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    377: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000010000000001000000011111000000000000000000000000000000000000000000000000001000100000000011111100000001011111100011001000001010000000000111000001111111111100011110000000000011010000011100000000000000011111000010000000111111111111111111101110100111111110111000101111111100000000000000000000000000000000000100000001011111111000000000000000000000000000000000011111100100100000110000000101000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    378: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111000000000000001110000000001000000010111000000000000000000000000000000000000000000000000000000000000000010111110000000011111101101010000001100000000001110000010111111111001011100000000001111110001111110010000000000001111000000000000111110110111111010000000000001111110010000111110111100000000000000000000000000000000000000000000111111100000000000000000000000000000000000011111100000100000011000000000000000000000000000000001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    379: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000100000000110100000011111100000000000000000000000000000000000000000000000000000000000010001111101000000010111110110011000001100000000011110000011111111110001111000000000000111111000111100000000000000111110000000000000111111111110111110000000000011111111000000111111110000000000000000000000000000000000000000000001111110100000000100000000000000000000000000011111000001000000001010000000000000000000000000000001111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    380: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000000101000100000001000000011111000000000000000000000000000000001000000000000000000000000000000000011110100000001111110111001100010110000000001100100011111010110101110001001000011111111101111110000000000000011110100000000000101111111111111111000000000000111111100000011111111000000010000000000000000010000000000000000010111111010000000000000000000000000000000000011111100000110000001100000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    381: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010000000000001100001000100001000011111110000000000000000000000000000000000000000000000000000000000000000001111101000000111110111100100001010000000111100010011111111110001111000000000011111011110111100000010000010111110000010000000110111111111110111100000000000011011110001111111100000000000000100000000000001000000000000000011011111000000000000000000000000000000000000011011000000010000001010000010000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    382: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000110000000001111001000000000000000000000000000000000000000000000000000000000000000001111110100000101111111001000001101000000011100000111111111000111000000000001011111111111111100000000001111111111100000000000111110111111110110000000000000011111111000111111010000000000000000000000000000000000000000000111111100000000000000000000000000000000000000011111100000100000000110000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    383: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010000000000010000000001000000000011111110100000000000000000000000000000000000000000000000000000000000010000011111100001111111111101100011100000001111000000011111111100111100000000000111111111111111000000000010111111111110000000000111111111110100011100000000000000111111011111101000000000000000000000000000000000000000000001111111010001000000000000000000000000000000000111111000000110000000010000000000000000000000000000001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    384: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000100000000000011111010101000100000000000000000000000000000000000000000000000000000000011111111000011111110100100000100000000111100001111111111001111100000000001111111101111110110000000111110111111111101000000011111111011110011110100000000001111011111101100000000000000000000000000000000000000000000101111111000000000000000000000000000000000000000011111000000101000000001000000000000000000000000000001111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    385: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111110000000000010000000000010000000000000111110000000000000000000000000000000000000000000000000000000000000000000111111000011111111100110001110000011011000001011111111010111000000000011111111111111111000000010111111101111111111010101111111111111100010100000000000000011111111110100000000000000000000000000000000000000000000010111101000000000000000000000000000000000000000111111100000010000000100100000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    386: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000010111111000001111111100100000100100001110000001110110110111111100000000110111111101111111100010111111111110001111011111111111111100001100001010000000000000001111111100000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000111110010001010000000010000001000010000000000000000001111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    387: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000011111000001000000000000000000000000000000000000000000000000000000000011110100011111111110100011100000011011000001011111110011111000000100011111101011101111101011111111111100001111111111111011101100011100000000000000000000010110111010000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    388: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000011111100000000000000000000000000000001000000000000111110000000000000000000000000000000000000000000000000000000000000111111000000011111110110000110001011110000001111111110111011110000001111111111111111111111111111111111100011101111111111111110000001100000000000000000000001111111100000000000000000000000000000000000000000000111111111000000000000000000000000000000000000100001111111000000000000000000010000000000000000000000000001011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    389: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000100000000000011110000000000000000000000000000000000000000000000000000000000000001111100001011111110110000010001010011000001111111100011101101000001111111111011111111111111111110101000001110011011111101000000001100000000000000000000000011111000000000000000000000000000000000000000010000011111100000000000000000000000000000000000000000000011111000000100000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    390: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000100000000000000000000000000000000000000101111010000000000000000000000000000000000000000000000000000000000000101111010000101110110111000010001111000000011111111100111111110100111111111010101111011111111101011110000011100001101011101000000001100000000000000000000000001111100000000000000000000000000000000000000000111111011100000000000000000000000000000000000000000001101101000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    391: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000011111100000011111111010001000011110110000001111111100011111111001011011011111011111101111111110001110001011000000000011100000000001100000000000000000000000011111100000000000000000000000000000000010000000011111110000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000010000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    392: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000010000000111110000000000000000000000000000000000000000000000000000000000000011111111000001111111111000000001110100000011111110100111111111110111111110111111111010010110100000100000011110000000001100000000001101000000000000000000000000111110000000000000000000000000000000000000001111111110100000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    393: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010111000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000011111111010000111111111100000001111010100001011111000011111111111111101011010111111000001111000011110000011001000000011110000000001100100000000000000000000010111110010000000000000000000000000000000000110110111110000010000000000000000000000000000000000000010111111000000000000000000000000000000000000000000000001101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    394: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111000000000000000000000000000000000000000000010111100000000000000000000000000000000000000000000000000000000000000110111111000010111111111000000001101100000111111111000111111111111111110101111111111000011111000011000000011000000000011100000000001100000000000000000000000001111110000000000000000000000000000000001011011111111000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    395: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000000000001011111111110000011111111100000001110100000001111111000111011111111111110011011011110000001100000011100000111000000001011001000010001100000000000000000000000001111110000000000000000000000000000000001111111111111110010000000000000000000000000000000000000000000111101000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    396: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000111100010000000000000000000000000000000000000000000000000000000000111111111101000101110111111000011111100000011111111000111111011111011110011111111111000011110010011000000011100000000001100000000000110000000000000000000000000111100000000000000000000000000000001011011100011111110000000000000000000000000000000000000000000000111110000000000010000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    397: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000000000000000000000000000000000000000001111100001000000000000000000000000000000000000000000000000000100000111111111111000001111111100000001111100000011101111000011111110111111110001111111100000011110000011100000010000000000101000000000010100000000000000000000000010111110000000000001000000000100000101111101000001111110000000000000000000000000000000000000000000010111101000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    398: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000011111101101111000000111111111000001111000000001111111001111111111110111110111111110100100011000000110001001011000000000000000000000000100000000000000000000000001111110000000000000000100000000000111111110000111111110000000000000000000000000000000000000000000001111110100000000000000000000000000000000000000000001000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    399: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000010111111011111100000111111110000001111100000011111110000111111101110011000011111111000000111100000111000000111000000000000000000000000000000000000000000000000001111110000000000000000000000000111111111000000011111010000000000000000000000000000000000000000000000111111010000000000000000000000000000000000000000000001110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    400: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010010000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000011111111101011110000101111111100001101000000011111111000111110111011011100111011101000001011000000101000000011000000000000000000000000000000000000000000000000000111111001000000000000000000000111111111000000111111100000000000000000000000000000000000000000000010111111011110000000000000000000000000000000000000000001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    401: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011011111100111111000010111111100001111000000001111110000111111101110011000011111110000000111100000111000000011000000000000000000000000000000000000000000000000011011110000000000000000000000001111101111000010111111110000000000000000000000000000000000000000000001011111111010100000000000000000000000000000000000000001111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    402: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000010000111100000000000000000000000000000000000000000000000000000000000111101111111011111000000111111110001111100000101110111000111101110110011001111111010000000110000000100000000101000000000000000000000000000000000000000000000000001111110000000000000000000101101111111000000001101111000000000000000000000000000000000000000000000001111111111111101000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    403: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010000000000000000000000000000000000000010000000111110000000000000000000000000000000000000000000000000000000001011000111110111011000001011111100001111000000111111110000111101111011011011111111000000000111000011110000000110000000000000000000000000000010000000000000000000011111101000000000000000101111111110101100000011111110000000000000000000000000000000000000000000000000111111101011111000010000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    404: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000001011100000000000000000000000000000000000000000000000000000000001111100111111110110110000101111111000111100000001111111000001110100110011011111101100000000101000000110000000101000000000000000000000000000000000000000000000000001111110000000000000010110111111101010000000101111111000010000000000000000000000000000000000000000000111111110101111111000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    405: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000010000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000010000000001110110011111111001010000001011111100101100000011111111000011110111011011110111110000000000110000001111000000011000000000000000000000000000000000000000001000000000111110000000000000011011111111110110000000111111110000000100000000000000000000000000000000000000000011011010000100110100000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    406: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111010100000000000000000000000000000000000000000100000111100000000000000000000000000000000000000000000000000000000010111010111111111100101000000111101101111100000001111101000001110001111011111111110000000000010000001100000000001000000000000000000000000000000000000000000000000011111100000000000000001001111100111010000010111111010000000000000000000000000000000000000000000000001011111101001110011010000100000000000000000000000000001111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    407: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000011111000111110000001000000000000000000000000000000000000000000001000111101111111111110010100000000001111101111000000011111111000001110000101111111111110000000000000000010100000000100000000000000000000000000000000000000000000000000011110110000000000001010010110110010000001001111101000000000000000000000000000000000000000000000000000111111101100010010101000000001000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    408: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111101000000000000000000000000000000000000000011110110111010100000000000000000000000000000000000000000000000000000111000111111011111000101100000010111110111100000000101101000010111010111111111101111000000000000000001110000000000000000000000000000000000000000000000000000000000010111100000000000000001011111101101000000111111111000000000000000000000000000000000000000000000000000011111100010001001000010000000000100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    409: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000010000000000000000000000000101111011111011110010000010000000000000000000000000000000000000000000001011100111101101111100100010000000011111111110000001001111000000110001111111110100100000000000000001001010000000010001000000000000000000000000000000000000000000000011111110000000000000101111101010100000000111110100000000000000000000000000000000000000000000000000000001111110010001001010000100000000000000000000000000000101101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    410: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000000000000100000000000000000000011111000111111111100000000010000000000000000000000000000000000000000001111000111100111111000110010000000001111111100000000001111000000111011111111110001110000000000000000001000000000000000000000000000000000000000000000000000000000000011111000000000000000101011101010000000111111111000000000000000000000000000000000000000000000000000000011111101001000100101000010000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    411: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000001000000000000000000000000000000111100010011111111111000000000000000000000000000000000000000000000000111101110011100011111100001101000000000101111110000000100111000000111101110111000000110010000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000111001000000010111111110000000000000001000000000000000000000000000000000000000001111110000001001000100010000000000010000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    412: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000001101100000000011111111111000000000000000000000000000000000000000000010011011101111000001111110010010000000000010111111000000000101000000011111111110100000101000000000000000000100000000000000000000000000000000000000000000000000000000000011111000000000000000001100010100010000111111101001000000000000000000000000000000000000000000000010001000111111000000010000000000101000000000000000000000000011101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    413: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000100010001001110000000000001101111101101000010000000000000000000000000000000101011101001111111000000101100001001000000000000101111010000000111100001011111111110000000110000000000000000000010000000000000000000000000000000000000000000000000000000000011011100000000000000000001010000000111111011110000000000000000000000000000000000000000000000000000000000011011000000001100100000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    414: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000111100000000000001111111111110000000000000000000000000000000000010111101111001111010000011111110001010100000000000010111000000000011000001111101110001010100111000000000000000000000000000000000000000000000000000000000000000000000001000000111100000000000000000000001101000001111011111111000000000000000000000000000000000000000000000000000000001011111100000000000000000101000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    415: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000001011010000000000001100111111111110000000000000000000000000000100000111010111100111100000001111010000000101000000000001111000000000011100111111111100111111011110000000000000000000000000000000000000000000000000000000000000000000000000000001011111000000000000000000001000000010111111100111100010000000000000000000000000000000000000000000000000000011111000000000000000010000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    416: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111000000000000001000000000000101111000000000000000110011010111111010000000000000000000000000000000101000101010111010000000111101000000100000000000001111100000000001101011011110101010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000011000000111111110100011111000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    417: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000010101111111110100011110000001000000001100111101111111110100000000000000000000000000000111000011011111000000000111110000000001000100000000110100000000001111111111110000110000100000000000000000000000000000000000001000000000000000000000000000000000000000010001111010000000000000000010000000001111111110000010110000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    418: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000111111111111111111111111010000000000000001110010101111111111100010000000100000000000000000001100111111100000000000111110000000000100000100000111000000000011111111111001001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000010000000000000000000111111111110001011111000000000000000000000000000000000000000000000000000000000111101000000000000000000000000000000000000000000111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    419: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110110000001011011010101111111111100000000000000001000011000110011111110000000000000000000000000000010111111100000000000000111111000000010000000000000111100100010101111111101000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000100000000100001011111111100101111111110000000000000000000000000000000000000000000000000000001011110100000000000000000000000000001000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    420: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110100000000000000000000001010100000000000100000110011001101011111111100000000000000000000000000000111011010000001000000011101000000000000000000000011010000011111111111100000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000010000000000000000000001111101111110111110101101000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    421: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110100000000000001000000000000000000000000000001110101001110001101111111000000000000000000000000000000100000000000000000011111100000000000000000000001100001111111110110100000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000001111111101111111010001110100010000000000000000000000000000000000000000000000000001110110000000000000000000000000000000000000000110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    422: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000001100011000110111100111111000000000000000000000000000000000000000000000000011111000000000000000000000001111110111111111000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000010111100000000000000000000000000111111111101111110000001111000000000000000000000000000000000000000000000000000000001111010001000000000000001000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    423: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111101000000000000000000000000000000000000010000100110001101001000111111110000000000000000000000000000000100000000000000101111000000000000000000000000111111111111110100001101000010110000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000001111111110011111010100000011110000000010000000000000000000000000000000000000000000001111110000000000000000100000100000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    424: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000100101000000001010011000110011100111011101000000000000000000000000000000001000000000000011101100000000000000000000001111111111111000000000110100000111000000000000000000000000000000000000000000000000000000000000000000000000000010111101000000000000000000000000000111011111000111100000010111100000000000000000000000000000000000000000000000000000000011111000000000000000000001011000010000000000101111000100000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    425: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000010111100000000000001001010101000010111111100000000000000000000000000000000000000000000011111110000000000000000000110101111110110100000001111110000101000000000000000000000000000000000000000000000000000000000000000000000100001001111101000000000000000000000000001111101100000011100000011111110000000000000000000000000000000000000000000000000000000111111000000000000000000101101100000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    426: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011110000000000000000000000000000011011100000000100111001100111000110011111110010000000000000000000000000000000000000000001111000000000000000001010111111101111000000000001110111000111000000000000000000000000000000000000000000000000000000000000000000000000001111111100010000000000000000000000001111111100001011100001111111110000000000000000000000000000000000000000000000000000000011111000000000000000001111111110000000000000011111100001000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    427: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000111101110000000000010000110001100000000111010000000000000000000000000000000001000000000011111110001000000001000111111111111110010000001001100101110011000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000001011111111000000011110011011011111000000000000000000000000000000000000000000000000000000111011000000000000000110111101111001000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    428: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100010000000000000000000000000011001010000000000011000100011000010000011111000000010000000000000000000000100001000000001111110000000000000011111111111111000000001000001110010101011000000000000000000000000000000000000000000000000000000000000000000000011011111101000000000000000000000000000001111111000000101110011101010110001000000000000000000000000000000000000000000000000000011111100000010000101111100001011110010010100001110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    429: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110100000000000000000000000000000011101110000000000001000110101000000100011111111010000000000000000000000110111101010000001111100000000100101111111111111010000000101100000110000011101000000000000000000000000000000000000000000000000000000000000000000000001111110100000000000000000000000100000001111111000000001111011110001110000000000000000000000000000000000000000000000000000100011111000000000010011110100000101101111111111101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    430: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000001011111010000000000000000000111000000000011111111101010010000000010001011011111111010100001110110000000000111111111111011000000000011110001110000000100000000000000000000000000000000000000000000000000000000000000100000001111111110000000000000000000000000000000110111100000000000111111000000111000000000000000000000000000000000000000000000000000000101111000000001011111010000000010111111111110101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    431: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000010000000111111000000000000000001100001100000001111111111111101000001000000010111111111101111011011011110000000111111101111111100000000000001110100111000000000000010000000000000000000000000000000000000000000000000000010000000101111101100001000000000000000000000000000011111110000000000111111100001110000000000000000000000000000000000000000000000000000000111111000000101111101000000000000110101001111110111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    432: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010110000000000000000000010001110000001110100000000000010000000011000000010111111111111111111110101001011111111011111111111111111110000011111111111110100000000100000000111000011000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000011111010000000001011111100000111000000000000000000000000000000000000000000000000000000011111001011111110100000000000000000100000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    433: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000010000000000000000011000000000010000000000000000000000001000001111110111111111111111011111111111111111111111111111111111111001101111111111110100000000000001000011100111100000000000000000000000000000000000000000000000000000000000000000000001001111111111111000000000100000000000000000001011111010000000000001111100011110000000000000000000000000000000000000000000000000000001011111000111111000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    434: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000100000000000000000000000000000000000000011111111000101111111111111111111111111100010110111111111111111111111110111110100000000000010110000001110010000000010000000000000000000000000000000000000000100000000000100000000000011111111111111000000000000000000000000000000111111100000000000101011100101111000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    435: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001111100000000000000000000000000000000000000000100000000000000000000001111111000000000001111111111111111111101001000000101011111111110111111111110100000000000000000101000010101111100000000000000000000000000000000000000000010000000000000000000000000000111111101111111100100000000000000000000000001011111000000000000000111111111110000000000000000000000000000000000000000000000000000001111011111111011000000000000000000000000000000000011111110001000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    436: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010000000000000000000000000000000000000000001000000000000000000111111101010000000000000111111111111110100000000000000010011111111111111111101000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000001110111111111111100000000000000000000000000001111111000000000000000001111111100000001000000000000000000000000000000000000000000000010111111111110101100000000000000000000000000000000101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    437: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000100000010000000010101111100000000000000100000001001010010000000000000000001001101111111101010000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111110110111110000000000000000000000000101111101000000000000000000110110100000000000000000000000000000000000000000000000001000001111110110111011010000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    438: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111000000000100000000000000000000000000000000000000000000000101011111110000000000000000000000100000001000000000000000000000111111111011110000000000000001000100100000000000000100000000000000000000000000100000000000000000000000000000000000000000000011111111111110011111000000000001000000000000111111110100000000000000000010110000000000000000000000000000000000000000000000000000000110111111111111011000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    439: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000101000001010011111111001000000000000000000000000000000000000000000000000011101111011100001000000000000000000000000000000000000000000000000000000000000000000010010110000000000000000000000000000000001111110111111100111111100000000100000001000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111110100011101100000000000000000000000000000000001011111100000100000000000000000000000000000000000000000000000000000000000000000000000000  ;
    440: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111111010111111111110100000000000000000000000000000000000000000000000101101111101100010000000000000000000000000000000000000000000010000000000000100001000010101111011101000000000000000000000000000001111111001111110001111010000000000000000010011101111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111011011000000000000000000000000000000000000000111101000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    441: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000001111111111111111111010000000100000000000000000000000000000000000000000011111110101000000000000000000000000000000000000000000000000000000000000000000000001011011011101110000000000000000000000000000001111111111111110001111101000000000000000001111110111110000000000000000000000000000000000000000000000000000000000000000000000000000001011111110110011011100100000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    442: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000001111000111111111100010000000000000010000000000000000000000000000000000111111110010000000000000000010000000000000000000000000000000000000000000000000000001101001000000100111000000000000000000000000001011111110101111100000111110000000000000000101111111111000000100000000000000000000010000000000000000000000000000000000000000000000000001111111100111011011000000000000000000000000000000000000100111111000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    443: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000001111100111101000010000000000000000000000000000000000000000000000000111111110101000000000000000001000000000000000000000000000000000000000000000000001101100000000000000000000100000000000000000000000000111010110111011110000111111000000000000101011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111010110010101100000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000  ; 
    444: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000010000000010111101101110100000000000000000000000000000000000000000000000010011011111110000000000000000000000000000000000000000000000000000000000000000000010111010001000000000100000010000000000000000000000000000111111000101111010000011111100000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111011011100000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000  ; 
    445: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001011110000001000000000000000000000000000000000011011101111110000000000000000000000000000000000000000000000000001011111010000000000000000000000000000000000000000000000000000000000000000000000001011100000000000000000000000100010000000000000000010000111100000111011110000101111100000010001011110111111110001000000000000000000000000000000000000000000000000000000000000000000000000000101111111100011011010100000000000000000000000000000010101000011111110001000000000000000000000000000000000000000000000000000000000000000000000000  ;
    446: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000010001100000000000000010000000000000000011111011111100000000000000000000000000000000000000000000000010111111111100100000000000000000000000000000000000000000000000000000000000000000101111010000000010001000000000000000000001000000000000000011111101000011011010000011011100000000001011111110111110000000000000000000000000000000000000000000000000000000000000000000000000000000011011111100110011011000000000000000000000000000000011111100001111101000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    447: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100001111010100000000000000000000000100001111111111111000000100000000000000000000001000000000000000101101111111000000000000000000000000000000000000000000000000000000000100000000000000110111000000000000010100000100000000000000000000000000000001111100000001101110000011111110000000000000111111110110000000000000000000000000000000000000000000000000000000000000000000000000000000111111111101011011001100010000000000000000000000001011101111000111110000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    448: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010111111110000000000000000000000000000000111111101111000000010010000000000000000010111010010001011011111111101000000000000000000000000000000000000000000000000000000000000000000000101011000000000101101001110011010101000000000000000000000000010111000000010011101000001111100000000000000000111111101000001000000000000000000000000100000000000000000000000000000000000000000000000111110111100110001011010000000000000000000100000000111000111101011111000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    449: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001111011111111110000000000000000000000000010101110111111111000001110000000000000000000011111101000100111111111101000000000000000000000000000000000000000000000000000000000000000000000000111110000000010111110110111111111111101000000000000000000000011110000000000101110000010111110000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111101100010001001100000000000000000000000000000101000001100011111100000000000000000000000000000000000000000000000000000000000000000000000000  ;
    450: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111000111110000000000000000000000010111111111010111010010000110000100000000000000011111111111111111111110101000000000000000000000000000000000000000000000000000000000000000010000101100000000011111111111011001011111111111110000010010000000000011110000000000110110000001111110000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000001000010111111111100110000000000000000000000000000000000000110000101100011111100000000000000000000000000000000000000000000000000000000000000000000000000  ;
    451: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101101011110001000000000000000111111111111111111111100000001111000000000000010001111111111111111111111011110100000000000000000000000000000000000000000000000000000000000000000010110110000011101111011111111101011111111111111101000000000000000001000000000000001010000001111110000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111100010000000100000000000000000000000000000111000011110001111110000000000000000000000000000000000000000000000000000000000000000000000000  ;
    452: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000111101000000000000000011011111111101111011111010000000111100000000000000000110111111110111111010111101000000000000000000000000000000000000000000000000100000000000000001010100000010101111010000111111100000101111111111110000000000000000010100000000000000100000001011101000000000000000000010111111100100000000000000000000000000000000000000000000000000000000000000000000011111111111100110000000000000000000000000000000000000011111011100000111111010000000000000000000000000000000000000000000000000000000000000000000000  ;
    453: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100001111110000010000000000011111110111111111111111000000001101000000000000000000111101111111111101011010100000000000000000000000000000000000000000000000000000000000000000001010100000011111111000000111111100000000001011111110100000000010000000000000000000000010000001111110000000000000000000001011111110000001000000000000000000000000000000000000000000000000000010000000000011111101101110010000000000000000000000000000000000000001111111100000111111000000000000000000000000000000000000000000000000000000000000000000000000  ;
    454: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000111110000000000000011111011111111101111111111000000001111100000000000000000111101111111010101111100000000000000000000000000000000000000000000000000000000000000000000010100000011111111000000000011111110000000000001101111100000000010000001001000000000000000000000111110000000000000000000000011111110100000000100000000000000000000000000000000000000000000000000000000001111111111110100010000000000000000000000000000000000000100111010100000011111100000000000000000000000000000000000000000000000000000000000000000000000  ;
    455: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000011010101111101111110111110000000001111000000000000000001111110111111101011010000000000000000000000000000000000000000000000000000000001000100000101101000011111111100100000000011111100000000000110111111111000001101000101110000000000000000000001111101000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001001011111111111100000000000000001000000000000000000000100000000000000000010111110000000000000000000000000000000000000000000000000000000000000000000000  ;
    456: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000111110000000000010111100001111101011101110111000000001111110000000000000001111111111000010111110100000000000000000000000000000000000000000000000000000001111000001010000000101111110000000000011101111110000001000011111111110100000000000111101000000000000000000001111100000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000011111101110110110001000000000000000000000000000000000000000000000000000001111101000000000000000000000000000000000000000000000000000000000000000000000  ;
    457: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010000000000001101000000111101111110111100000000000111100000000000000000111111001010101101010001000100000000000000000000000000000000000000000000000101101110101101000111111111101000000000001100111010001100000011111111111110000100010111111010001010000000000001111110000000000000000000000000010111111000000000000000000000000000000000000000000000000000000000000000001101111111111010000000000000000000000000000000000000000000000000000000000011110100000000000000000000000000000000000000000000000000000000000000000000  ;
    458: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000011100000000011110111111111110000000011110110000000000000011111111000010111111010000000000000000000000000000000000000000000000000000000010101111101000001011111101000000010001110111011100101111000001111101111010000000011100110000101110010001001010111000001000000000001000000000011110111000000000000000000000000000000000000000000000000000000000000001111111111110111100000000000100000000000000000000000000000000000000000000000101111000000000000000000000000000000000000000000000000000000000000000000000  ;
    459: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000010000110000000000111111001011111000000000000111100000000000000001011100001011101110000000000000000000000000000000000000000000000000000100000011000001010001111111101110000000000000101011111110011111000000011111111110000000111010111000111011100000000011111100000000000000100010000000001011111100000000000000000000000000000000000000000000000000000000000000111111110111101100000000000000000000000000000000000000000000000001000000000011111100000000000000000000000000000000000000000000000000000000000000000000  ;
    460: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000010111000000000011111100111011100000100001111110000000000010001111010111110111000000000000000000000000000000000000000000000000001000000010111100000000010011111111110000000000000110001111000000100110000011111111111100000000000011000110111100000000111111000000000000000000001101000000111111110000000000000000000000000000000000000000000000000000000000001111111111010111010000000000000000000000000000000000000000000000000010000010111111000000000000000000000000000000000000000000000000000000000000000000000  ;
    461: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100010010010100000000000000001010111110100000000001111010000000000000101111111010111010000000000000000000000000000000000000000000000100000000000011011100000001011111111100111000000000000010000111000011110100000001110111110100000000000011111010011100111100111111000000000000000000000100000000011111110000000000000000000000000000000000000000000000000000000000101111111011101111100000000000000000000000000000100000000000000000000000000001011111100000000000000000000000000000000000000000000000000000000000000000000  ;
    462: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111011111111100000000000000000011111111000000000001111100000000000000011111111011101000000000000000000000000000000000000000000000000000000000011101000010000011111101101000111000000000011100000000000000111100000000111111111110000000000011111000011010111111111010000000000000000000000011000000111101110000000000000000000000000000000000000000000000000000010000111111101010110111100000000000000000000000000000000000000000000000000000010111111110100000000000000000000000000000000000000000000000000000000000000000000  ;
    463: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000100000000000000111111110000000000001011110000000000000001111111110000000100000000000000000000000000000000000000000000000000001010100001000010101111111010001110100100100001101000000000001111000000001111111111101000001000001111000011011111111011101000000000000000000000001100000011111101000010000000000000000000000000000000000000000000000000001011110110111011101100010000000000001000100000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000  ;
    464: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111101110101111000000000000000001011111111000000000001111100000000000000001011111101000000000000000000000000000000000000000000000100000000000001101000000000001111110110000001011101111000000100000000000000010100000000011111111111000000000000000000011111101111111100000000001000000000000000011100101111111000000000000000000000000000000000000000000000000000000001111111100001111111010000000000100100000000000000000000000000000000000000101111111000000000000000000000000000000000000000000000000000000000000000000000000  ;
    465: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110101111100000000001000000011101111110000000000001111110000000000000011111100000000000000000000000000000000000000000000000000000000000000100100000000001111111111000000001111111111101001100000000000010000001000000101111111111100000000000000100011111100111111000000000000000000000000000001000001111111000000000000000000000000000000000000000000000000000000111111111000000010101000001010111111111111010000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000  ;
    466: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001011110000000000000001011111111101000000000001111110000000000000001101100000000000000000000000000000000000000000000000000000000000101010000000000111111111000000000011111111011110011100000000000000000000000000010111010100000000100000000000011100011111110000000000000000000000000000001110101111110000000000000000000000000000000000000000000000000000001111101100000000000100100001111111111111111111101000000000000001000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    467: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000001000111110101110000000000001111101000000000000011111100000000000000000000000000000000100000000000000000000000010101000000000010101111100000000000101011000000011001100000000000000000000000000001111100000010100000010000000000110011111010000000000000000000000000000000111011111011000000000000000000000000000000000000000000000000000111011111100000000000010011111111111111111111111110000001000001000000000000001111111010000000000000000000000000000000000000000000000000000000000000000000000000  ;
    468: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000011111110111100000000000000011110000000000000000111100000000000000000000000000000000000000000000000000000100011100000001000111111110100000000000111101000000011010110000000000000000000000000001111100000001111111000000000000000111111000000010000000000000100000010000011111111110000000000000000000000000000000000000000000000010000111111110100000000000101111111111110111110101111111111000000000000000000000001011101000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    469: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001111100000000000000011111001011100000000000001111111000000000000001111110000000000000000000000000000000000001000000000000000001101000000000101111111110000000000000010011100000011001100100000000000000000000000000111110010001111110100000000000001011111000000000000000000000000000000000001101111111000000000000000000000000000000000000000000000000011011111111000101000111111111111111111111110000011111111100000000000000000000001111111000001000000000000000000000000000000000000000000000000000000000000000000000  ;
    470: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000001111010000111100000000000000111100000000000000000111100000000000000000000000000000000000000000000000000001101100000000000111111100000100000000001111010000000011011100000000000000000000100000010111010000001111011110000000000001111000000100000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111101100001111101111111101010111111100000000111111111000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    471: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110100000000000010111110000111110000000000001110111000000000000001111110000000000000000000000000000000000000000000000000010110010000000111111111101000000000100000110111000010111001100000000000000000000000001000111100000000011111111100000001011110000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000011111111111111111111111111101010101111101001000000000111111110000000000000000001111110100000000000000000000000000000000000000000000000000000000000000000000000000  ;
    472: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000100000011111100000111000000000000000111111000000000000001011111000100000000000000000000000000000000001000000001010100000000011011111010000000000000000000010111000000001101000000000000000000000000000000111110000000001111111111101001111100100000000000000000000000000000000000000010111110000000000000000000000000000000000000000000000000001011101111111111111111101010100000011110100000000000001011101100000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000  ;         
    473: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000010011111000000111100000000000000111111000000000000000101111000000000000000000000000000000000000000000010101010000000001011111111101000000000000000001111111000000111101100000000000000000000000000000011100000000000010110110111111101000000000000000000000000000000000000000001011011111000000000000000000000000000000000000000000000000000000111111111111111111100000000000111110000000000000001011111101000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000  ;
    474: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111110010000000001011101000000111110000000000000011111000000010000000111111000000000000000000000000000000000000000000001010000000001001111111100000000000000000000000011101000000010110100000000000000000000000000000111110000000000000011011101111100100000000000000000000000000000000000000000111111100010000000000000000000000000000000000000000000000000000111101011010011111010000000000011110000000000000000001011110100000000000010111110100000000000000000000000000000000000000000000000000000000000000000000000000  ;
    475: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110111000000000001111110000000111100000000000000111111000100000000000011011000001000000000000000000000000000000000010110100000010001111111110101000000000000000000000001100000000011111000000000000000000000000000000111110000100000000001011111100000000000000000000000000000000000000000000000001110110000000000000000000000000000000000000000000000000000000111100000000011101000000000000111100000000000000000000101111110000100000001111111000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    476: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000011111100000000111100000000000000011011100000000000000011111100000000100000000000000000000000000001001010000000000011111111101000000000000000000000000000000000000000110000000100000000000000000000000011100000000000000000000111111000000000000000000000000000000000000000000000011111110000000010000000000000000000000000000000000000000000000101110000000001111000000000000011100000000000000000000000111101000000010000110111100000000000000000000000000000000000000000000000000000000000000000000000000  ;
    477: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000001111100100000011110000000000000011111100000000000000001111110000000000000000000000000000000000001111000000100011101111110100000000000000000000000000000000000000100010000000000000000000000000000000011110000000101000000000001100000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000001111010000000011100000000000000011010000000000000000000000011111100000000000111101000000000000000000000000000000000000000000000000000000000000000000000000000  ;
    478: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000111010100000001011000000000000000101111000000000000000001111110000000000000000000000000000100010110101000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000010111110000111110100000000001110000000000000000000000000000000000000000000000001110100000000000000000000000000000000000000000000000000000001111100000001011100000000000000011100000000000000000000000001111110000000000111111000100000000000000000000000000000000000000000000000000000000000000000000000  ;
    479: dataREG = 641'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000111111000000000111110000000000000011101110000000000000010111110000000000000000000000000010010011110000000000011111111010010000000000000000000000000000000000000000000000000000000000000000000000000000011100000110111110000000001010000000000000000000000000000000000000000000000011111100000000000000100000000000000000000000000000000000000001111010010000111000000000000000111000000000000000000000000001111111000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000  ;
     default: dataREG=0;
     endcase 
     end               
    assign W_o = wREG;
    assign H_o = hREG;
    assign data_o = dataREG;
    endmodule

