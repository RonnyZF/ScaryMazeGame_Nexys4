`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Ronny Zarate Ferreto
// 
// Create Date: 07.09.2017 23:01:31
// Design Name: 
// Module Name: Sincronizador_VGA
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Sincronizador_VGA(
    input wire clk, reset,
    output wire hsync, vsync, video_on, p_tick,
    output wire [9:0] pixel_x, pixel_y
   );

   // constant declaration
   // VGA 640-by-480 sync parameters
   localparam HD = 640; // horizontal display area
   localparam HF = 48 ; // h. front (left) border
   localparam HB = 16 ; // h. back (right) border
   localparam HR = 96 ; // h. retrace
   localparam VD = 480; // vertical display area
   localparam VF = 10;  // v. front (top) border
   localparam VB = 33;  // v. back (bottom) border
   localparam VR = 2;   // v. retrace

   // mod-2 counter
   reg mod2_reg;
   wire mod2_next;
   reg mod2_reg2;
   wire mod2_next2;

   // sync counters
   reg [9:0] h_count_reg, h_count_next;
   reg [9:0] v_count_reg, v_count_next;
   // output buffer
   reg v_sync_reg, h_sync_reg;
   wire v_sync_next, h_sync_next;
   // status signal
   wire h_end, v_end, pixel_tick;

   // registers
   always @(posedge clk, posedge reset)
      if (reset)
         begin
            mod2_reg <= 1'b0;

         end
      else
         begin
            mod2_reg <= mod2_next;

         end
   // mod-2 circuit to generate 25 MHz enable tick
   assign mod2_next = ~mod2_reg;
  // assign pixel_tick = mod2_reg;
   
    always @(posedge clk, posedge reset)
      if (reset)
       begin
          mod2_reg2 <=1'b0;
          v_sync_reg <= 1'b0;
          h_sync_reg <= 1'b0;
       end
    else
        if (mod2_reg)
       begin
          mod2_reg2 <= mod2_next2;
          v_sync_reg <= v_sync_next;
          h_sync_reg <= h_sync_next;
       end
    
   assign mod2_next2 = ~mod2_reg2;
   assign pixel_tick = mod2_reg2;
   
   // status signals
   // end of horizontal counter (799)
  assign h_end = (h_count_reg==(HD+HF+HB+HR-1));
   // end of vertical counter (524)
   assign v_end = (v_count_reg==(VD+VF+VB+VR-1));

   // next-state logic of mod-800 horizontal sync counter
   always @(posedge pixel_tick+1)
         if (reset)
            h_count_reg <= 0;
         else if (h_end)
             h_count_reg <= 0;
         else
            begin
            h_count_reg <= h_count_reg + 1;
            //h_count_reg <= h_count_next;
            end
     
   // next-state logic of mod-525 vertical sync counter
   always @(posedge pixel_tick+1)
      if (reset)
        v_count_reg <= 0;
      else if (h_end)
         if (v_end)
            v_count_reg <= 0;
         else
            begin
            v_count_reg <= v_count_reg + 1;
            //v_count_reg <= v_count_next;

            end
      else
         v_count_reg <= v_count_reg;

   // horizontal and vertical sync, buffered to avoid glitch
   // h_sync_next asserted between 656 and 751
   assign h_sync_next = ~(h_count_reg>=(HD+HB) && h_count_reg<=(HD+HB+HR-1));
   // vh_sync_next asserted between 490 and 491
   assign v_sync_next = ~(v_count_reg>=(VD+VB) && v_count_reg<=(VD+VB+VR-1));

   // video on/off
   assign video_on = (h_count_reg<HD) && (v_count_reg<VD);

   // output
 
   assign hsync = h_sync_reg;
   assign vsync = v_sync_reg;
   assign pixel_x = h_count_reg;
   assign pixel_y = v_count_reg;
   assign p_tick = pixel_tick;

endmodule
